// ------------------------------------------------------------------
//  Design Unit:    aes256_encrypt_ecb_core
// ------------------------------------------------------------------


module aes256_encrypt_ecb_core (
  clk, rst, ctx_key_triosy_lz, ctx_enckey_triosy_lz, ctx_deckey_triosy_lz, k_triosy_lz,
      buf_rsc_zout, buf_rsc_lzout, buf_rsc_zin, buf_triosy_lz, ctx_key_rsci_data_in_d,
      ctx_key_rsci_addr_rd_d, ctx_key_rsci_addr_wr_d, ctx_key_rsci_re_d, ctx_key_rsci_we_d,
      ctx_key_rsci_data_out_d, ctx_enckey_rsci_addr_rd_d, ctx_enckey_rsci_addr_wr_d,
      ctx_enckey_rsci_re_d, ctx_enckey_rsci_we_d, ctx_enckey_rsci_data_out_d, ctx_deckey_rsci_data_in_d,
      ctx_deckey_rsci_addr_rd_d, ctx_deckey_rsci_addr_wr_d, ctx_deckey_rsci_re_d,
      ctx_deckey_rsci_we_d, ctx_deckey_rsci_data_out_d, k_rsci_addr_rd_d, k_rsci_re_d,
      k_rsci_data_out_d, aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_addr, aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out,
      aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_en
);
  input clk;
  input rst;
  output ctx_key_triosy_lz;
  output ctx_enckey_triosy_lz;
  output ctx_deckey_triosy_lz;
  output k_triosy_lz;
  output [127:0] buf_rsc_zout;
  output buf_rsc_lzout;
  input [127:0] buf_rsc_zin;
  output buf_triosy_lz;
  output [7:0] ctx_key_rsci_data_in_d;
  output [4:0] ctx_key_rsci_addr_rd_d;
  output [4:0] ctx_key_rsci_addr_wr_d;
  output ctx_key_rsci_re_d;
  output ctx_key_rsci_we_d;
  input [7:0] ctx_key_rsci_data_out_d;
  output [4:0] ctx_enckey_rsci_addr_rd_d;
  output [4:0] ctx_enckey_rsci_addr_wr_d;
  output ctx_enckey_rsci_re_d;
  output ctx_enckey_rsci_we_d;
  input [7:0] ctx_enckey_rsci_data_out_d;
  output [7:0] ctx_deckey_rsci_data_in_d;
  output [4:0] ctx_deckey_rsci_addr_rd_d;
  output [4:0] ctx_deckey_rsci_addr_wr_d;
  output ctx_deckey_rsci_re_d;
  output ctx_deckey_rsci_we_d;
  input [7:0] ctx_deckey_rsci_data_out_d;
  output [4:0] k_rsci_addr_rd_d;
  output k_rsci_re_d;
  input [7:0] k_rsci_data_out_d;
  output [7:0] aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_addr;
  reg [7:0] aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_addr;
  input [7:0] aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out;
  output aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_en;

  assign cpkey_mux1h_159_nl = MUX1HOT_v_3_7_2((cpkey_cpkey_xor_1_cmx_sva_1[7:5]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[127:125]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[7:5]),
      mix_mix_xor_7_cmx_7_5_sva_1, (buf_rsci_din[127:125]), (ctx_key_rsci_data_in_d_mx0w1[7:5]),
      (buf_rsci_din[95:93]), {and_dcpl_231 , and_dcpl_232 , and_dcpl_235 , and_dcpl_206
      , and_dcpl_219 , and_dcpl_236 , and_dcpl_92});
  assign cpkey_mux1h_157_nl = MUX1HOT_v_2_7_2((cpkey_cpkey_xor_1_cmx_sva_1[4:3]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[124:123]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[4:3]),
      mix_mix_xor_7_cmx_4_3_sva_1, (buf_rsci_din[124:123]), (ctx_key_rsci_data_in_d_mx0w1[4:3]),
      (buf_rsci_din[92:91]), {and_dcpl_231 , and_dcpl_232 , and_dcpl_235 , and_dcpl_206
      , and_dcpl_219 , and_dcpl_236 , and_dcpl_92});
  assign cpkey_mux1h_155_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[2]), (addkey_1_io_read_buf_rsc_sdt_1_sva[122]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[2]), mix_mix_xor_7_cmx_2_sva_1,
      (buf_rsci_din[122]), (ctx_key_rsci_data_in_d_mx0w1[2]), (buf_rsci_din[90]),
      {and_dcpl_231 , and_dcpl_232 , and_dcpl_235 , and_dcpl_206 , and_dcpl_219 ,
      and_dcpl_236 , and_dcpl_92});
  assign cpkey_mux1h_153_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[1]), (addkey_1_io_read_buf_rsc_sdt_1_sva[121]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[1]), mix_mix_xor_7_cmx_1_sva_1,
      (buf_rsci_din[121]), (ctx_key_rsci_data_in_d_mx0w1[1]), (buf_rsci_din[89]),
      {and_dcpl_231 , and_dcpl_232 , and_dcpl_235 , and_dcpl_206 , and_dcpl_219 ,
      and_dcpl_236 , and_dcpl_92});
  assign cpkey_mux1h_151_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[0]), (addkey_1_io_read_buf_rsc_sdt_1_sva[120]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[0]), mix_mix_xor_7_cmx_0_sva_1,
      (buf_rsci_din[120]), (ctx_key_rsci_data_in_d_mx0w1[0]), (buf_rsci_din[88]),
      {and_dcpl_231 , and_dcpl_232 , and_dcpl_235 , and_dcpl_206 , and_dcpl_219 ,
      and_dcpl_236 , and_dcpl_92});
  assign cpkey_mux1h_149_nl = MUX1HOT_v_3_7_2((cpkey_cpkey_xor_1_cmx_sva_1[7:5]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[119:117]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[7:5]),
      mix_mix_xor_5_cmx_7_5_sva_1, (buf_rsci_din[119:117]), (ctx_key_rsci_data_in_d_mx0w1[7:5]),
      (buf_rsci_din[55:53]), {and_dcpl_223 , and_dcpl_224 , and_dcpl_227 , and_dcpl_206
      , and_dcpl_219 , and_dcpl_228 , and_dcpl_92});
  assign cpkey_mux1h_147_nl = MUX1HOT_v_2_7_2((cpkey_cpkey_xor_1_cmx_sva_1[4:3]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[116:115]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[4:3]),
      mix_mix_xor_5_cmx_4_3_sva_1, (buf_rsci_din[116:115]), (ctx_key_rsci_data_in_d_mx0w1[4:3]),
      (buf_rsci_din[52:51]), {and_dcpl_223 , and_dcpl_224 , and_dcpl_227 , and_dcpl_206
      , and_dcpl_219 , and_dcpl_228 , and_dcpl_92});
  assign cpkey_mux1h_145_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[2]), (addkey_1_io_read_buf_rsc_sdt_1_sva[114]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[2]), mix_mix_xor_5_cmx_2_sva_1,
      (buf_rsci_din[114]), (ctx_key_rsci_data_in_d_mx0w1[2]), (buf_rsci_din[50]),
      {and_dcpl_223 , and_dcpl_224 , and_dcpl_227 , and_dcpl_206 , and_dcpl_219 ,
      and_dcpl_228 , and_dcpl_92});
  assign cpkey_mux1h_143_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[1]), (addkey_1_io_read_buf_rsc_sdt_1_sva[113]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[1]), mix_mix_xor_5_cmx_1_sva_1,
      (buf_rsci_din[113]), (ctx_key_rsci_data_in_d_mx0w1[1]), (buf_rsci_din[49]),
      {and_dcpl_223 , and_dcpl_224 , and_dcpl_227 , and_dcpl_206 , and_dcpl_219 ,
      and_dcpl_228 , and_dcpl_92});
  assign cpkey_mux1h_141_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[0]), (addkey_1_io_read_buf_rsc_sdt_1_sva[112]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[0]), mix_mix_xor_5_cmx_0_sva_1,
      (buf_rsci_din[112]), (ctx_key_rsci_data_in_d_mx0w1[0]), (buf_rsci_din[48]),
      {and_dcpl_223 , and_dcpl_224 , and_dcpl_227 , and_dcpl_206 , and_dcpl_219 ,
      and_dcpl_228 , and_dcpl_92});
  assign cpkey_mux1h_139_nl = MUX1HOT_v_3_7_2((cpkey_cpkey_xor_1_cmx_sva_1[7:5]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[111:109]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[7:5]),
      mix_mix_xor_3_cmx_7_5_sva_1, (buf_rsci_din[111:109]), (ctx_key_rsci_data_in_d_mx0w1[7:5]),
      (buf_rsci_din[15:13]), {and_dcpl_213 , and_dcpl_214 , and_dcpl_217 , and_dcpl_206
      , and_dcpl_219 , and_dcpl_220 , and_dcpl_92});
  assign cpkey_mux1h_137_nl = MUX1HOT_v_2_7_2((cpkey_cpkey_xor_1_cmx_sva_1[4:3]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[108:107]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[4:3]),
      mix_mix_xor_3_cmx_4_3_sva_1, (buf_rsci_din[108:107]), (ctx_key_rsci_data_in_d_mx0w1[4:3]),
      (buf_rsci_din[12:11]), {and_dcpl_213 , and_dcpl_214 , and_dcpl_217 , and_dcpl_206
      , and_dcpl_219 , and_dcpl_220 , and_dcpl_92});
  assign cpkey_mux1h_135_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[2]), (addkey_1_io_read_buf_rsc_sdt_1_sva[106]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[2]), mix_mix_xor_3_cmx_2_sva_1,
      (buf_rsci_din[106]), (ctx_key_rsci_data_in_d_mx0w1[2]), (buf_rsci_din[10]),
      {and_dcpl_213 , and_dcpl_214 , and_dcpl_217 , and_dcpl_206 , and_dcpl_219 ,
      and_dcpl_220 , and_dcpl_92});
  assign cpkey_mux1h_133_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[1]), (addkey_1_io_read_buf_rsc_sdt_1_sva[105]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[1]), mix_mix_xor_3_cmx_1_sva_1,
      (buf_rsci_din[105]), (ctx_key_rsci_data_in_d_mx0w1[1]), (buf_rsci_din[9]),
      {and_dcpl_213 , and_dcpl_214 , and_dcpl_217 , and_dcpl_206 , and_dcpl_219 ,
      and_dcpl_220 , and_dcpl_92});
  assign cpkey_mux1h_131_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[0]), (addkey_1_io_read_buf_rsc_sdt_1_sva[104]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[0]), mix_mix_xor_3_cmx_0_sva_1,
      (buf_rsci_din[104]), (ctx_key_rsci_data_in_d_mx0w1[0]), (buf_rsci_din[8]),
      {and_dcpl_213 , and_dcpl_214 , and_dcpl_217 , and_dcpl_206 , and_dcpl_219 ,
      and_dcpl_220 , and_dcpl_92});
  assign cpkey_mux1h_129_nl = MUX1HOT_v_3_6_2((cpkey_cpkey_xor_1_cmx_sva_1[7:5]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[103:101]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[7:5]),
      mix_mix_xor_1_cmx_7_5_sva_1, (ctx_key_rsci_data_in_d_mx0w1[7:5]), (buf_rsci_din[103:101]),
      {and_dcpl_200 , not_tmp_151 , and_dcpl_203 , and_dcpl_206 , and_dcpl_209 ,
      and_dcpl_210});
  assign cpkey_mux1h_127_nl = MUX1HOT_v_2_6_2((cpkey_cpkey_xor_1_cmx_sva_1[4:3]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[100:99]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[4:3]),
      mix_mix_xor_1_cmx_4_3_sva_1, (ctx_key_rsci_data_in_d_mx0w1[4:3]), (buf_rsci_din[100:99]),
      {and_dcpl_200 , not_tmp_151 , and_dcpl_203 , and_dcpl_206 , and_dcpl_209 ,
      and_dcpl_210});
  assign cpkey_mux1h_125_nl = MUX1HOT_s_1_6_2((cpkey_cpkey_xor_1_cmx_sva_1[2]), (addkey_1_io_read_buf_rsc_sdt_1_sva[98]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[2]), mix_mix_xor_1_cmx_2_sva_1,
      (ctx_key_rsci_data_in_d_mx0w1[2]), (buf_rsci_din[98]), {and_dcpl_200 , not_tmp_151
      , and_dcpl_203 , and_dcpl_206 , and_dcpl_209 , and_dcpl_210});
  assign cpkey_mux1h_123_nl = MUX1HOT_s_1_6_2((cpkey_cpkey_xor_1_cmx_sva_1[1]), (addkey_1_io_read_buf_rsc_sdt_1_sva[97]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[1]), mix_mix_xor_1_cmx_1_sva_1,
      (ctx_key_rsci_data_in_d_mx0w1[1]), (buf_rsci_din[97]), {and_dcpl_200 , not_tmp_151
      , and_dcpl_203 , and_dcpl_206 , and_dcpl_209 , and_dcpl_210});
  assign cpkey_mux1h_121_nl = MUX1HOT_s_1_6_2((cpkey_cpkey_xor_1_cmx_sva_1[0]), (addkey_1_io_read_buf_rsc_sdt_1_sva[96]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[0]), mix_mix_xor_1_cmx_0_sva_1,
      (ctx_key_rsci_data_in_d_mx0w1[0]), (buf_rsci_din[96]), {and_dcpl_200 , not_tmp_151
      , and_dcpl_203 , and_dcpl_206 , and_dcpl_209 , and_dcpl_210});
  assign cpkey_mux1h_119_nl = MUX1HOT_v_3_7_2((cpkey_cpkey_xor_1_cmx_sva_1[7:5]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[95:93]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[7:5]),
      mix_mix_xor_7_cmx_7_5_sva_1, (buf_rsci_din[95:93]), (ctx_key_rsci_data_in_d_mx0w1[7:5]),
      (buf_rsci_din[63:61]), {and_dcpl_192 , and_dcpl_193 , and_dcpl_196 , and_dcpl_165
      , and_dcpl_177 , and_dcpl_197 , and_dcpl_92});
  assign cpkey_mux1h_117_nl = MUX1HOT_v_2_7_2((cpkey_cpkey_xor_1_cmx_sva_1[4:3]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[92:91]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[4:3]),
      mix_mix_xor_7_cmx_4_3_sva_1, (buf_rsci_din[92:91]), (ctx_key_rsci_data_in_d_mx0w1[4:3]),
      (buf_rsci_din[60:59]), {and_dcpl_192 , and_dcpl_193 , and_dcpl_196 , and_dcpl_165
      , and_dcpl_177 , and_dcpl_197 , and_dcpl_92});
  assign cpkey_mux1h_115_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[2]), (addkey_1_io_read_buf_rsc_sdt_1_sva[90]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[2]), mix_mix_xor_7_cmx_2_sva_1,
      (buf_rsci_din[90]), (ctx_key_rsci_data_in_d_mx0w1[2]), (buf_rsci_din[58]),
      {and_dcpl_192 , and_dcpl_193 , and_dcpl_196 , and_dcpl_165 , and_dcpl_177 ,
      and_dcpl_197 , and_dcpl_92});
  assign cpkey_mux1h_113_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[1]), (addkey_1_io_read_buf_rsc_sdt_1_sva[89]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[1]), mix_mix_xor_7_cmx_1_sva_1,
      (buf_rsci_din[89]), (ctx_key_rsci_data_in_d_mx0w1[1]), (buf_rsci_din[57]),
      {and_dcpl_192 , and_dcpl_193 , and_dcpl_196 , and_dcpl_165 , and_dcpl_177 ,
      and_dcpl_197 , and_dcpl_92});
  assign cpkey_mux1h_111_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[0]), (addkey_1_io_read_buf_rsc_sdt_1_sva[88]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[0]), mix_mix_xor_7_cmx_0_sva_1,
      (buf_rsci_din[88]), (ctx_key_rsci_data_in_d_mx0w1[0]), (buf_rsci_din[56]),
      {and_dcpl_192 , and_dcpl_193 , and_dcpl_196 , and_dcpl_165 , and_dcpl_177 ,
      and_dcpl_197 , and_dcpl_92});
  assign cpkey_mux1h_109_nl = MUX1HOT_v_3_7_2((cpkey_cpkey_xor_1_cmx_sva_1[7:5]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[87:85]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[7:5]),
      mix_mix_xor_5_cmx_7_5_sva_1, (buf_rsci_din[87:85]), (ctx_key_rsci_data_in_d_mx0w1[7:5]),
      (buf_rsci_din[23:21]), {and_dcpl_184 , (~ mux_174_itm) , and_dcpl_187 , and_dcpl_165
      , and_dcpl_177 , and_dcpl_189 , and_dcpl_92});
  assign cpkey_mux1h_107_nl = MUX1HOT_v_2_7_2((cpkey_cpkey_xor_1_cmx_sva_1[4:3]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[84:83]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[4:3]),
      mix_mix_xor_5_cmx_4_3_sva_1, (buf_rsci_din[84:83]), (ctx_key_rsci_data_in_d_mx0w1[4:3]),
      (buf_rsci_din[20:19]), {and_dcpl_184 , (~ mux_174_itm) , and_dcpl_187 , and_dcpl_165
      , and_dcpl_177 , and_dcpl_189 , and_dcpl_92});
  assign cpkey_mux1h_105_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[2]), (addkey_1_io_read_buf_rsc_sdt_1_sva[82]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[2]), mix_mix_xor_5_cmx_2_sva_1,
      (buf_rsci_din[82]), (ctx_key_rsci_data_in_d_mx0w1[2]), (buf_rsci_din[18]),
      {and_dcpl_184 , (~ mux_174_itm) , and_dcpl_187 , and_dcpl_165 , and_dcpl_177
      , and_dcpl_189 , and_dcpl_92});
  assign cpkey_mux1h_103_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[1]), (addkey_1_io_read_buf_rsc_sdt_1_sva[81]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[1]), mix_mix_xor_5_cmx_1_sva_1,
      (buf_rsci_din[81]), (ctx_key_rsci_data_in_d_mx0w1[1]), (buf_rsci_din[17]),
      {and_dcpl_184 , (~ mux_174_itm) , and_dcpl_187 , and_dcpl_165 , and_dcpl_177
      , and_dcpl_189 , and_dcpl_92});
  assign cpkey_mux1h_101_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[0]), (addkey_1_io_read_buf_rsc_sdt_1_sva[80]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[0]), mix_mix_xor_5_cmx_0_sva_1,
      (buf_rsci_din[80]), (ctx_key_rsci_data_in_d_mx0w1[0]), (buf_rsci_din[16]),
      {and_dcpl_184 , (~ mux_174_itm) , and_dcpl_187 , and_dcpl_165 , and_dcpl_177
      , and_dcpl_189 , and_dcpl_92});
  assign cpkey_mux1h_99_nl = MUX1HOT_v_3_7_2((cpkey_cpkey_xor_1_cmx_sva_1[7:5]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[79:77]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[7:5]),
      mix_mix_xor_3_cmx_7_5_sva_1, (buf_rsci_din[79:77]), (ctx_key_rsci_data_in_d_mx0w1[7:5]),
      (buf_rsci_din[111:109]), {and_dcpl_172 , not_tmp_142 , and_dcpl_175 , and_dcpl_165
      , and_dcpl_177 , and_dcpl_180 , and_dcpl_92});
  assign cpkey_mux1h_97_nl = MUX1HOT_v_2_7_2((cpkey_cpkey_xor_1_cmx_sva_1[4:3]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[76:75]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[4:3]),
      mix_mix_xor_3_cmx_4_3_sva_1, (buf_rsci_din[76:75]), (ctx_key_rsci_data_in_d_mx0w1[4:3]),
      (buf_rsci_din[108:107]), {and_dcpl_172 , not_tmp_142 , and_dcpl_175 , and_dcpl_165
      , and_dcpl_177 , and_dcpl_180 , and_dcpl_92});
  assign cpkey_mux1h_95_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[2]), (addkey_1_io_read_buf_rsc_sdt_1_sva[74]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[2]), mix_mix_xor_3_cmx_2_sva_1,
      (buf_rsci_din[74]), (ctx_key_rsci_data_in_d_mx0w1[2]), (buf_rsci_din[106]),
      {and_dcpl_172 , not_tmp_142 , and_dcpl_175 , and_dcpl_165 , and_dcpl_177 ,
      and_dcpl_180 , and_dcpl_92});
  assign cpkey_mux1h_93_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[1]), (addkey_1_io_read_buf_rsc_sdt_1_sva[73]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[1]), mix_mix_xor_3_cmx_1_sva_1,
      (buf_rsci_din[73]), (ctx_key_rsci_data_in_d_mx0w1[1]), (buf_rsci_din[105]),
      {and_dcpl_172 , not_tmp_142 , and_dcpl_175 , and_dcpl_165 , and_dcpl_177 ,
      and_dcpl_180 , and_dcpl_92});
  assign cpkey_mux1h_91_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[0]), (addkey_1_io_read_buf_rsc_sdt_1_sva[72]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[0]), mix_mix_xor_3_cmx_0_sva_1,
      (buf_rsci_din[72]), (ctx_key_rsci_data_in_d_mx0w1[0]), (buf_rsci_din[104]),
      {and_dcpl_172 , not_tmp_142 , and_dcpl_175 , and_dcpl_165 , and_dcpl_177 ,
      and_dcpl_180 , and_dcpl_92});
  assign cpkey_mux1h_89_nl = MUX1HOT_v_3_6_2((cpkey_cpkey_xor_1_cmx_sva_1[7:5]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[71:69]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[7:5]),
      mix_mix_xor_1_cmx_7_5_sva_1, (ctx_key_rsci_data_in_d_mx0w1[7:5]), (buf_rsci_din[71:69]),
      {and_dcpl_158 , not_tmp_137 , and_dcpl_162 , and_dcpl_165 , and_dcpl_168 ,
      and_dcpl_169});
  assign cpkey_mux1h_87_nl = MUX1HOT_v_2_6_2((cpkey_cpkey_xor_1_cmx_sva_1[4:3]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[68:67]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[4:3]),
      mix_mix_xor_1_cmx_4_3_sva_1, (ctx_key_rsci_data_in_d_mx0w1[4:3]), (buf_rsci_din[68:67]),
      {and_dcpl_158 , not_tmp_137 , and_dcpl_162 , and_dcpl_165 , and_dcpl_168 ,
      and_dcpl_169});
  assign cpkey_mux1h_85_nl = MUX1HOT_s_1_6_2((cpkey_cpkey_xor_1_cmx_sva_1[2]), (addkey_1_io_read_buf_rsc_sdt_1_sva[66]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[2]), mix_mix_xor_1_cmx_2_sva_1,
      (ctx_key_rsci_data_in_d_mx0w1[2]), (buf_rsci_din[66]), {and_dcpl_158 , not_tmp_137
      , and_dcpl_162 , and_dcpl_165 , and_dcpl_168 , and_dcpl_169});
  assign cpkey_mux1h_83_nl = MUX1HOT_s_1_6_2((cpkey_cpkey_xor_1_cmx_sva_1[1]), (addkey_1_io_read_buf_rsc_sdt_1_sva[65]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[1]), mix_mix_xor_1_cmx_1_sva_1,
      (ctx_key_rsci_data_in_d_mx0w1[1]), (buf_rsci_din[65]), {and_dcpl_158 , not_tmp_137
      , and_dcpl_162 , and_dcpl_165 , and_dcpl_168 , and_dcpl_169});
  assign cpkey_mux1h_81_nl = MUX1HOT_s_1_6_2((cpkey_cpkey_xor_1_cmx_sva_1[0]), (addkey_1_io_read_buf_rsc_sdt_1_sva[64]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[0]), mix_mix_xor_1_cmx_0_sva_1,
      (ctx_key_rsci_data_in_d_mx0w1[0]), (buf_rsci_din[64]), {and_dcpl_158 , not_tmp_137
      , and_dcpl_162 , and_dcpl_165 , and_dcpl_168 , and_dcpl_169});
  assign cpkey_mux1h_79_nl = MUX1HOT_v_3_7_2((cpkey_cpkey_xor_1_cmx_sva_1[7:5]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[63:61]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[7:5]),
      mix_mix_xor_7_cmx_7_5_sva_1, (buf_rsci_din[63:61]), (ctx_key_rsci_data_in_d_mx0w1[7:5]),
      (buf_rsci_din[31:29]), {and_dcpl_149 , and_dcpl_150 , and_dcpl_153 , and_dcpl_125
      , and_dcpl_136 , and_dcpl_154 , and_dcpl_92});
  assign cpkey_mux1h_77_nl = MUX1HOT_v_2_7_2((cpkey_cpkey_xor_1_cmx_sva_1[4:3]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[60:59]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[4:3]),
      mix_mix_xor_7_cmx_4_3_sva_1, (buf_rsci_din[60:59]), (ctx_key_rsci_data_in_d_mx0w1[4:3]),
      (buf_rsci_din[28:27]), {and_dcpl_149 , and_dcpl_150 , and_dcpl_153 , and_dcpl_125
      , and_dcpl_136 , and_dcpl_154 , and_dcpl_92});
  assign cpkey_mux1h_75_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[2]), (addkey_1_io_read_buf_rsc_sdt_1_sva[58]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[2]), mix_mix_xor_7_cmx_2_sva_1,
      (buf_rsci_din[58]), (ctx_key_rsci_data_in_d_mx0w1[2]), (buf_rsci_din[26]),
      {and_dcpl_149 , and_dcpl_150 , and_dcpl_153 , and_dcpl_125 , and_dcpl_136 ,
      and_dcpl_154 , and_dcpl_92});
  assign cpkey_mux1h_73_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[1]), (addkey_1_io_read_buf_rsc_sdt_1_sva[57]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[1]), mix_mix_xor_7_cmx_1_sva_1,
      (buf_rsci_din[57]), (ctx_key_rsci_data_in_d_mx0w1[1]), (buf_rsci_din[25]),
      {and_dcpl_149 , and_dcpl_150 , and_dcpl_153 , and_dcpl_125 , and_dcpl_136 ,
      and_dcpl_154 , and_dcpl_92});
  assign cpkey_mux1h_71_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[0]), (addkey_1_io_read_buf_rsc_sdt_1_sva[56]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[0]), mix_mix_xor_7_cmx_0_sva_1,
      (buf_rsci_din[56]), (ctx_key_rsci_data_in_d_mx0w1[0]), (buf_rsci_din[24]),
      {and_dcpl_149 , and_dcpl_150 , and_dcpl_153 , and_dcpl_125 , and_dcpl_136 ,
      and_dcpl_154 , and_dcpl_92});
  assign cpkey_mux1h_69_nl = MUX1HOT_v_3_7_2((cpkey_cpkey_xor_1_cmx_sva_1[7:5]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[55:53]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[7:5]),
      mix_mix_xor_5_cmx_7_5_sva_1, (buf_rsci_din[55:53]), (ctx_key_rsci_data_in_d_mx0w1[7:5]),
      (buf_rsci_din[119:117]), {and_dcpl_141 , not_tmp_128 , and_dcpl_144 , and_dcpl_125
      , and_dcpl_136 , and_dcpl_146 , and_dcpl_92});
  assign cpkey_mux1h_67_nl = MUX1HOT_v_2_7_2((cpkey_cpkey_xor_1_cmx_sva_1[4:3]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[52:51]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[4:3]),
      mix_mix_xor_5_cmx_4_3_sva_1, (buf_rsci_din[52:51]), (ctx_key_rsci_data_in_d_mx0w1[4:3]),
      (buf_rsci_din[116:115]), {and_dcpl_141 , not_tmp_128 , and_dcpl_144 , and_dcpl_125
      , and_dcpl_136 , and_dcpl_146 , and_dcpl_92});
  assign cpkey_mux1h_65_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[2]), (addkey_1_io_read_buf_rsc_sdt_1_sva[50]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[2]), mix_mix_xor_5_cmx_2_sva_1,
      (buf_rsci_din[50]), (ctx_key_rsci_data_in_d_mx0w1[2]), (buf_rsci_din[114]),
      {and_dcpl_141 , not_tmp_128 , and_dcpl_144 , and_dcpl_125 , and_dcpl_136 ,
      and_dcpl_146 , and_dcpl_92});
  assign cpkey_mux1h_63_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[1]), (addkey_1_io_read_buf_rsc_sdt_1_sva[49]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[1]), mix_mix_xor_5_cmx_1_sva_1,
      (buf_rsci_din[49]), (ctx_key_rsci_data_in_d_mx0w1[1]), (buf_rsci_din[113]),
      {and_dcpl_141 , not_tmp_128 , and_dcpl_144 , and_dcpl_125 , and_dcpl_136 ,
      and_dcpl_146 , and_dcpl_92});
  assign cpkey_mux1h_61_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[0]), (addkey_1_io_read_buf_rsc_sdt_1_sva[48]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[0]), mix_mix_xor_5_cmx_0_sva_1,
      (buf_rsci_din[48]), (ctx_key_rsci_data_in_d_mx0w1[0]), (buf_rsci_din[112]),
      {and_dcpl_141 , not_tmp_128 , and_dcpl_144 , and_dcpl_125 , and_dcpl_136 ,
      and_dcpl_146 , and_dcpl_92});
  assign cpkey_mux1h_59_nl = MUX1HOT_v_3_7_2((cpkey_cpkey_xor_1_cmx_sva_1[7:5]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[47:45]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[7:5]),
      mix_mix_xor_3_cmx_7_5_sva_1, (buf_rsci_din[47:45]), (ctx_key_rsci_data_in_d_mx0w1[7:5]),
      (buf_rsci_din[79:77]), {and_dcpl_132 , (~ mux_146_itm) , and_dcpl_134 , and_dcpl_125
      , and_dcpl_136 , and_dcpl_138 , and_dcpl_92});
  assign cpkey_mux1h_57_nl = MUX1HOT_v_2_7_2((cpkey_cpkey_xor_1_cmx_sva_1[4:3]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[44:43]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[4:3]),
      mix_mix_xor_3_cmx_4_3_sva_1, (buf_rsci_din[44:43]), (ctx_key_rsci_data_in_d_mx0w1[4:3]),
      (buf_rsci_din[76:75]), {and_dcpl_132 , (~ mux_146_itm) , and_dcpl_134 , and_dcpl_125
      , and_dcpl_136 , and_dcpl_138 , and_dcpl_92});
  assign cpkey_mux1h_55_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[2]), (addkey_1_io_read_buf_rsc_sdt_1_sva[42]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[2]), mix_mix_xor_3_cmx_2_sva_1,
      (buf_rsci_din[42]), (ctx_key_rsci_data_in_d_mx0w1[2]), (buf_rsci_din[74]),
      {and_dcpl_132 , (~ mux_146_itm) , and_dcpl_134 , and_dcpl_125 , and_dcpl_136
      , and_dcpl_138 , and_dcpl_92});
  assign cpkey_mux1h_53_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[1]), (addkey_1_io_read_buf_rsc_sdt_1_sva[41]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[1]), mix_mix_xor_3_cmx_1_sva_1,
      (buf_rsci_din[41]), (ctx_key_rsci_data_in_d_mx0w1[1]), (buf_rsci_din[73]),
      {and_dcpl_132 , (~ mux_146_itm) , and_dcpl_134 , and_dcpl_125 , and_dcpl_136
      , and_dcpl_138 , and_dcpl_92});
  assign cpkey_mux1h_51_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[0]), (addkey_1_io_read_buf_rsc_sdt_1_sva[40]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[0]), mix_mix_xor_3_cmx_0_sva_1,
      (buf_rsci_din[40]), (ctx_key_rsci_data_in_d_mx0w1[0]), (buf_rsci_din[72]),
      {and_dcpl_132 , (~ mux_146_itm) , and_dcpl_134 , and_dcpl_125 , and_dcpl_136
      , and_dcpl_138 , and_dcpl_92});
  assign cpkey_mux1h_49_nl = MUX1HOT_v_3_6_2((cpkey_cpkey_xor_1_cmx_sva_1[7:5]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[39:37]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[7:5]),
      mix_mix_xor_1_cmx_7_5_sva_1, (ctx_key_rsci_data_in_d_mx0w1[7:5]), (buf_rsci_din[39:37]),
      {and_dcpl_118 , (~ mux_139_itm) , and_dcpl_122 , and_dcpl_125 , and_dcpl_129
      , and_dcpl_130});
  assign cpkey_mux1h_47_nl = MUX1HOT_v_2_6_2((cpkey_cpkey_xor_1_cmx_sva_1[4:3]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[36:35]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[4:3]),
      mix_mix_xor_1_cmx_4_3_sva_1, (ctx_key_rsci_data_in_d_mx0w1[4:3]), (buf_rsci_din[36:35]),
      {and_dcpl_118 , (~ mux_139_itm) , and_dcpl_122 , and_dcpl_125 , and_dcpl_129
      , and_dcpl_130});
  assign cpkey_mux1h_45_nl = MUX1HOT_s_1_6_2((cpkey_cpkey_xor_1_cmx_sva_1[2]), (addkey_1_io_read_buf_rsc_sdt_1_sva[34]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[2]), mix_mix_xor_1_cmx_2_sva_1,
      (ctx_key_rsci_data_in_d_mx0w1[2]), (buf_rsci_din[34]), {and_dcpl_118 , (~ mux_139_itm)
      , and_dcpl_122 , and_dcpl_125 , and_dcpl_129 , and_dcpl_130});
  assign cpkey_mux1h_43_nl = MUX1HOT_s_1_6_2((cpkey_cpkey_xor_1_cmx_sva_1[1]), (addkey_1_io_read_buf_rsc_sdt_1_sva[33]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[1]), mix_mix_xor_1_cmx_1_sva_1,
      (ctx_key_rsci_data_in_d_mx0w1[1]), (buf_rsci_din[33]), {and_dcpl_118 , (~ mux_139_itm)
      , and_dcpl_122 , and_dcpl_125 , and_dcpl_129 , and_dcpl_130});
  assign cpkey_mux1h_41_nl = MUX1HOT_s_1_6_2((cpkey_cpkey_xor_1_cmx_sva_1[0]), (addkey_1_io_read_buf_rsc_sdt_1_sva[32]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[0]), mix_mix_xor_1_cmx_0_sva_1,
      (ctx_key_rsci_data_in_d_mx0w1[0]), (buf_rsci_din[32]), {and_dcpl_118 , (~ mux_139_itm)
      , and_dcpl_122 , and_dcpl_125 , and_dcpl_129 , and_dcpl_130});
  assign cpkey_mux1h_39_nl = MUX1HOT_v_3_7_2((cpkey_cpkey_xor_1_cmx_sva_1[7:5]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[31:29]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[7:5]),
      (buf_rsci_din[31:29]), mix_mix_xor_7_cmx_7_5_sva_1, (ctx_key_rsci_data_in_d_mx0w1[7:5]),
      (buf_rsci_din[127:125]), {and_dcpl_108 , not_tmp_114 , and_dcpl_111 , and_dcpl_84
      , and_dcpl_61 , and_dcpl_114 , and_dcpl_92});
  assign cpkey_mux1h_37_nl = MUX1HOT_v_2_7_2((cpkey_cpkey_xor_1_cmx_sva_1[4:3]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[28:27]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[4:3]),
      (buf_rsci_din[28:27]), mix_mix_xor_7_cmx_4_3_sva_1, (ctx_key_rsci_data_in_d_mx0w1[4:3]),
      (buf_rsci_din[124:123]), {and_dcpl_108 , not_tmp_114 , and_dcpl_111 , and_dcpl_84
      , and_dcpl_61 , and_dcpl_114 , and_dcpl_92});
  assign cpkey_mux1h_35_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[2]), (addkey_1_io_read_buf_rsc_sdt_1_sva[26]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[2]), (buf_rsci_din[26]),
      mix_mix_xor_7_cmx_2_sva_1, (ctx_key_rsci_data_in_d_mx0w1[2]), (buf_rsci_din[122]),
      {and_dcpl_108 , not_tmp_114 , and_dcpl_111 , and_dcpl_84 , and_dcpl_61 , and_dcpl_114
      , and_dcpl_92});
  assign cpkey_mux1h_33_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[1]), (addkey_1_io_read_buf_rsc_sdt_1_sva[25]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[1]), (buf_rsci_din[25]),
      mix_mix_xor_7_cmx_1_sva_1, (ctx_key_rsci_data_in_d_mx0w1[1]), (buf_rsci_din[121]),
      {and_dcpl_108 , not_tmp_114 , and_dcpl_111 , and_dcpl_84 , and_dcpl_61 , and_dcpl_114
      , and_dcpl_92});
  assign cpkey_mux1h_31_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[0]), (addkey_1_io_read_buf_rsc_sdt_1_sva[24]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[0]), (buf_rsci_din[24]),
      mix_mix_xor_7_cmx_0_sva_1, (ctx_key_rsci_data_in_d_mx0w1[0]), (buf_rsci_din[120]),
      {and_dcpl_108 , not_tmp_114 , and_dcpl_111 , and_dcpl_84 , and_dcpl_61 , and_dcpl_114
      , and_dcpl_92});
  assign cpkey_mux1h_29_nl = MUX1HOT_v_3_7_2((cpkey_cpkey_xor_1_cmx_sva_1[7:5]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[23:21]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[7:5]),
      (buf_rsci_din[23:21]), mix_mix_xor_5_cmx_7_5_sva_1, (ctx_key_rsci_data_in_d_mx0w1[7:5]),
      (buf_rsci_din[87:85]), {and_dcpl_97 , (~ mux_128_itm) , and_dcpl_102 , and_dcpl_84
      , and_dcpl_61 , and_dcpl_106 , and_dcpl_92});
  assign cpkey_mux1h_27_nl = MUX1HOT_v_2_7_2((cpkey_cpkey_xor_1_cmx_sva_1[4:3]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[20:19]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[4:3]),
      (buf_rsci_din[20:19]), mix_mix_xor_5_cmx_4_3_sva_1, (ctx_key_rsci_data_in_d_mx0w1[4:3]),
      (buf_rsci_din[84:83]), {and_dcpl_97 , (~ mux_128_itm) , and_dcpl_102 , and_dcpl_84
      , and_dcpl_61 , and_dcpl_106 , and_dcpl_92});
  assign cpkey_mux1h_25_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[2]), (addkey_1_io_read_buf_rsc_sdt_1_sva[18]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[2]), (buf_rsci_din[18]),
      mix_mix_xor_5_cmx_2_sva_1, (ctx_key_rsci_data_in_d_mx0w1[2]), (buf_rsci_din[82]),
      {and_dcpl_97 , (~ mux_128_itm) , and_dcpl_102 , and_dcpl_84 , and_dcpl_61 ,
      and_dcpl_106 , and_dcpl_92});
  assign cpkey_mux1h_23_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[1]), (addkey_1_io_read_buf_rsc_sdt_1_sva[17]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[1]), (buf_rsci_din[17]),
      mix_mix_xor_5_cmx_1_sva_1, (ctx_key_rsci_data_in_d_mx0w1[1]), (buf_rsci_din[81]),
      {and_dcpl_97 , (~ mux_128_itm) , and_dcpl_102 , and_dcpl_84 , and_dcpl_61 ,
      and_dcpl_106 , and_dcpl_92});
  assign cpkey_mux1h_21_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[0]), (addkey_1_io_read_buf_rsc_sdt_1_sva[16]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[0]), (buf_rsci_din[16]),
      mix_mix_xor_5_cmx_0_sva_1, (ctx_key_rsci_data_in_d_mx0w1[0]), (buf_rsci_din[80]),
      {and_dcpl_97 , (~ mux_128_itm) , and_dcpl_102 , and_dcpl_84 , and_dcpl_61 ,
      and_dcpl_106 , and_dcpl_92});
  assign cpkey_mux1h_19_nl = MUX1HOT_v_3_7_2((cpkey_cpkey_xor_1_cmx_sva_1[7:5]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[15:13]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[7:5]),
      (buf_rsci_din[15:13]), mix_mix_xor_3_cmx_7_5_sva_1, (ctx_key_rsci_data_in_d_mx0w1[7:5]),
      (buf_rsci_din[47:45]), {and_dcpl_74 , (~ mux_121_itm) , and_dcpl_82 , and_dcpl_84
      , and_dcpl_61 , and_dcpl_89 , and_dcpl_92});
  assign cpkey_mux1h_17_nl = MUX1HOT_v_2_7_2((cpkey_cpkey_xor_1_cmx_sva_1[4:3]),
      (addkey_1_io_read_buf_rsc_sdt_1_sva[12:11]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[4:3]),
      (buf_rsci_din[12:11]), mix_mix_xor_3_cmx_4_3_sva_1, (ctx_key_rsci_data_in_d_mx0w1[4:3]),
      (buf_rsci_din[44:43]), {and_dcpl_74 , (~ mux_121_itm) , and_dcpl_82 , and_dcpl_84
      , and_dcpl_61 , and_dcpl_89 , and_dcpl_92});
  assign cpkey_mux1h_15_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[2]), (addkey_1_io_read_buf_rsc_sdt_1_sva[10]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[2]), (buf_rsci_din[10]),
      mix_mix_xor_3_cmx_2_sva_1, (ctx_key_rsci_data_in_d_mx0w1[2]), (buf_rsci_din[42]),
      {and_dcpl_74 , (~ mux_121_itm) , and_dcpl_82 , and_dcpl_84 , and_dcpl_61 ,
      and_dcpl_89 , and_dcpl_92});
  assign cpkey_mux1h_13_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[1]), (addkey_1_io_read_buf_rsc_sdt_1_sva[9]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[1]), (buf_rsci_din[9]),
      mix_mix_xor_3_cmx_1_sva_1, (ctx_key_rsci_data_in_d_mx0w1[1]), (buf_rsci_din[41]),
      {and_dcpl_74 , (~ mux_121_itm) , and_dcpl_82 , and_dcpl_84 , and_dcpl_61 ,
      and_dcpl_89 , and_dcpl_92});
  assign cpkey_mux1h_11_nl = MUX1HOT_s_1_7_2((cpkey_cpkey_xor_1_cmx_sva_1[0]), (addkey_1_io_read_buf_rsc_sdt_1_sva[8]),
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[0]), (buf_rsci_din[8]),
      mix_mix_xor_3_cmx_0_sva_1, (ctx_key_rsci_data_in_d_mx0w1[0]), (buf_rsci_din[40]),
      {and_dcpl_74 , (~ mux_121_itm) , and_dcpl_82 , and_dcpl_84 , and_dcpl_61 ,
      and_dcpl_89 , and_dcpl_92});
  assign cpkey_mux1h_9_nl = MUX1HOT_v_3_6_2((addkey_1_io_read_buf_rsc_sdt_1_sva[7:5]),
      (cpkey_cpkey_xor_1_cmx_sva_1[7:5]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[7:5]),
      mix_mix_xor_1_cmx_7_5_sva_1, (ctx_key_rsci_data_in_d_mx0w1[7:5]), (buf_rsci_din[7:5]),
      {not_tmp_81 , and_dcpl_48 , and_dcpl_53 , and_dcpl_61 , and_dcpl_63 , and_dcpl_66});
  assign cpkey_mux1h_7_nl = MUX1HOT_v_2_6_2((addkey_1_io_read_buf_rsc_sdt_1_sva[4:3]),
      (cpkey_cpkey_xor_1_cmx_sva_1[4:3]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[4:3]),
      mix_mix_xor_1_cmx_4_3_sva_1, (ctx_key_rsci_data_in_d_mx0w1[4:3]), (buf_rsci_din[4:3]),
      {not_tmp_81 , and_dcpl_48 , and_dcpl_53 , and_dcpl_61 , and_dcpl_63 , and_dcpl_66});
  assign cpkey_mux1h_5_nl = MUX1HOT_s_1_6_2((addkey_1_io_read_buf_rsc_sdt_1_sva[2]),
      (cpkey_cpkey_xor_1_cmx_sva_1[2]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[2]),
      mix_mix_xor_1_cmx_2_sva_1, (ctx_key_rsci_data_in_d_mx0w1[2]), (buf_rsci_din[2]),
      {not_tmp_81 , and_dcpl_48 , and_dcpl_53 , and_dcpl_61 , and_dcpl_63 , and_dcpl_66});
  assign cpkey_mux1h_3_nl = MUX1HOT_s_1_6_2((addkey_1_io_read_buf_rsc_sdt_1_sva[1]),
      (cpkey_cpkey_xor_1_cmx_sva_1[1]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[1]),
      mix_mix_xor_1_cmx_1_sva_1, (ctx_key_rsci_data_in_d_mx0w1[1]), (buf_rsci_din[1]),
      {not_tmp_81 , and_dcpl_48 , and_dcpl_53 , and_dcpl_61 , and_dcpl_63 , and_dcpl_66});
  assign cpkey_mux1h_1_nl = MUX1HOT_s_1_6_2((addkey_1_io_read_buf_rsc_sdt_1_sva[0]),
      (cpkey_cpkey_xor_1_cmx_sva_1[0]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[0]),
      mix_mix_xor_1_cmx_0_sva_1, (ctx_key_rsci_data_in_d_mx0w1[0]), (buf_rsci_din[0]),
      {not_tmp_81 , and_dcpl_48 , and_dcpl_53 , and_dcpl_61 , and_dcpl_63 , and_dcpl_66});
  assign nl_buf_rsci_dout = {cpkey_mux1h_159_nl , cpkey_mux1h_157_nl , cpkey_mux1h_155_nl
      , cpkey_mux1h_153_nl , cpkey_mux1h_151_nl , cpkey_mux1h_149_nl , cpkey_mux1h_147_nl
      , cpkey_mux1h_145_nl , cpkey_mux1h_143_nl , cpkey_mux1h_141_nl , cpkey_mux1h_139_nl
      , cpkey_mux1h_137_nl , cpkey_mux1h_135_nl , cpkey_mux1h_133_nl , cpkey_mux1h_131_nl
      , cpkey_mux1h_129_nl , cpkey_mux1h_127_nl , cpkey_mux1h_125_nl , cpkey_mux1h_123_nl
      , cpkey_mux1h_121_nl , cpkey_mux1h_119_nl , cpkey_mux1h_117_nl , cpkey_mux1h_115_nl
      , cpkey_mux1h_113_nl , cpkey_mux1h_111_nl , cpkey_mux1h_109_nl , cpkey_mux1h_107_nl
      , cpkey_mux1h_105_nl , cpkey_mux1h_103_nl , cpkey_mux1h_101_nl , cpkey_mux1h_99_nl
      , cpkey_mux1h_97_nl , cpkey_mux1h_95_nl , cpkey_mux1h_93_nl , cpkey_mux1h_91_nl
      , cpkey_mux1h_89_nl , cpkey_mux1h_87_nl , cpkey_mux1h_85_nl , cpkey_mux1h_83_nl
      , cpkey_mux1h_81_nl , cpkey_mux1h_79_nl , cpkey_mux1h_77_nl , cpkey_mux1h_75_nl
      , cpkey_mux1h_73_nl , cpkey_mux1h_71_nl , cpkey_mux1h_69_nl , cpkey_mux1h_67_nl
      , cpkey_mux1h_65_nl , cpkey_mux1h_63_nl , cpkey_mux1h_61_nl , cpkey_mux1h_59_nl
      , cpkey_mux1h_57_nl , cpkey_mux1h_55_nl , cpkey_mux1h_53_nl , cpkey_mux1h_51_nl
      , cpkey_mux1h_49_nl , cpkey_mux1h_47_nl , cpkey_mux1h_45_nl , cpkey_mux1h_43_nl
      , cpkey_mux1h_41_nl , cpkey_mux1h_39_nl , cpkey_mux1h_37_nl , cpkey_mux1h_35_nl
      , cpkey_mux1h_33_nl , cpkey_mux1h_31_nl , cpkey_mux1h_29_nl , cpkey_mux1h_27_nl
      , cpkey_mux1h_25_nl , cpkey_mux1h_23_nl , cpkey_mux1h_21_nl , cpkey_mux1h_19_nl
      , cpkey_mux1h_17_nl , cpkey_mux1h_15_nl , cpkey_mux1h_13_nl , cpkey_mux1h_11_nl
      , cpkey_mux1h_9_nl , cpkey_mux1h_7_nl , cpkey_mux1h_5_nl , cpkey_mux1h_3_nl
      , cpkey_mux1h_1_nl};
  wire  nl_aes256_encrypt_ecb_core_core_fsm_inst_ecb1_C_1_tr0;
  assign nl_aes256_encrypt_ecb_core_core_fsm_inst_ecb1_C_1_tr0 = z_out_1[5];
  wire  nl_aes256_encrypt_ecb_core_core_fsm_inst_exp1_C_9_tr0;
  assign nl_aes256_encrypt_ecb_core_core_fsm_inst_exp1_C_9_tr0 = z_out[2];
  wire  nl_aes256_encrypt_ecb_core_core_fsm_inst_exp2_C_9_tr0;
  assign nl_aes256_encrypt_ecb_core_core_fsm_inst_exp2_C_9_tr0 = z_out_1[3];
  wire  nl_aes256_encrypt_ecb_core_core_fsm_inst_mix_C_1_tr0;
  assign nl_aes256_encrypt_ecb_core_core_fsm_inst_mix_C_1_tr0 = (z_out[2]) & (~ (aes_addRoundKey_cpy_i_4_0_sva_1_3_0[0]));
  wire  nl_aes256_encrypt_ecb_core_core_fsm_inst_mix_C_1_tr1;
  assign nl_aes256_encrypt_ecb_core_core_fsm_inst_mix_C_1_tr1 = (z_out[2]) & (aes_addRoundKey_cpy_i_4_0_sva_1_3_0[0]);
  wire  nl_aes256_encrypt_ecb_core_core_fsm_inst_ecb3_C_10_tr0;
  assign nl_aes256_encrypt_ecb_core_core_fsm_inst_ecb3_C_10_tr0 = aes_addRoundKey_cpy_i_4_0_sva_1_3_0[0];
  wire  nl_aes256_encrypt_ecb_core_core_fsm_inst_exp1_1_C_9_tr0;
  assign nl_aes256_encrypt_ecb_core_core_fsm_inst_exp1_1_C_9_tr0 = z_out[2];
  wire  nl_aes256_encrypt_ecb_core_core_fsm_inst_ecb3_C_22_tr0;
  assign nl_aes256_encrypt_ecb_core_core_fsm_inst_ecb3_C_22_tr0 = aes_addRoundKey_cpy_i_4_0_sva_1_3_0[0];
  wire  nl_aes256_encrypt_ecb_core_core_fsm_inst_exp2_1_C_9_tr0;
  assign nl_aes256_encrypt_ecb_core_core_fsm_inst_exp2_1_C_9_tr0 = z_out_1[3];
  wire  nl_aes256_encrypt_ecb_core_core_fsm_inst_ecb3_C_23_tr0;
  assign nl_aes256_encrypt_ecb_core_core_fsm_inst_ecb3_C_23_tr0 = ~ (z_out_1[3]);
  wire  nl_aes256_encrypt_ecb_core_core_fsm_inst_exp1_2_C_9_tr0;
  assign nl_aes256_encrypt_ecb_core_core_fsm_inst_exp1_2_C_9_tr0 = z_out[2];
  wire  nl_aes256_encrypt_ecb_core_core_fsm_inst_exp2_2_C_9_tr0;
  assign nl_aes256_encrypt_ecb_core_core_fsm_inst_exp2_2_C_9_tr0 = z_out_1[3];
  aes256_encrypt_ecb_core_wait_dp aes256_encrypt_ecb_core_wait_dp_inst (
      .aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_en(aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_en),
      .aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_cgo(aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_cgo)
    );
  aes256_encrypt_ecb_core_core_fsm aes256_encrypt_ecb_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .ecb1_C_1_tr0(nl_aes256_encrypt_ecb_core_core_fsm_inst_ecb1_C_1_tr0),
      .ecb2_C_9_tr0(ecb2_ecb2_or_tmp),
      .exp1_C_9_tr0(nl_aes256_encrypt_ecb_core_core_fsm_inst_exp1_C_9_tr0),
      .ecb2_C_21_tr0(ecb2_ecb2_or_tmp),
      .exp2_C_9_tr0(nl_aes256_encrypt_ecb_core_core_fsm_inst_exp2_C_9_tr0),
      .ecb2_C_25_tr0(and_498_cse),
      .sub_C_0_tr0(and_dcpl_38),
      .mix_C_1_tr0(nl_aes256_encrypt_ecb_core_core_fsm_inst_mix_C_1_tr0),
      .mix_C_1_tr1(nl_aes256_encrypt_ecb_core_core_fsm_inst_mix_C_1_tr1),
      .addkey_C_0_tr0(and_dcpl_38),
      .ecb3_C_10_tr0(nl_aes256_encrypt_ecb_core_core_fsm_inst_ecb3_C_10_tr0),
      .exp1_1_C_9_tr0(nl_aes256_encrypt_ecb_core_core_fsm_inst_exp1_1_C_9_tr0),
      .ecb3_C_22_tr0(nl_aes256_encrypt_ecb_core_core_fsm_inst_ecb3_C_22_tr0),
      .exp2_1_C_9_tr0(nl_aes256_encrypt_ecb_core_core_fsm_inst_exp2_1_C_9_tr0),
      .addkey_1_C_0_tr0(and_dcpl_38),
      .ecb3_C_23_tr0(nl_aes256_encrypt_ecb_core_core_fsm_inst_ecb3_C_23_tr0),
      .sub_1_C_0_tr0(and_dcpl_38),
      .exp1_2_C_9_tr0(nl_aes256_encrypt_ecb_core_core_fsm_inst_exp1_2_C_9_tr0),
      .exp2_2_C_9_tr0(nl_aes256_encrypt_ecb_core_core_fsm_inst_exp2_2_C_9_tr0),
      .addkey_2_C_0_tr0(and_dcpl_38)
    );
  assign or_288_cse = (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1!=4'b0000) | addkey_1_nor_6_itm;
  assign or_290_cse = (fsm_output[1:0]!=2'b00);
  assign nand_99_cse = ~((fsm_output[4]) & (fsm_output[6]));
  assign nor_272_cse = ~((fsm_output[1:0]!=2'b00));
  assign nor_274_cse = ~((fsm_output[5]) | (fsm_output[0]));
  assign nor_279_cse = ~((fsm_output[4:3]!=2'b00));
  assign or_337_cse = (~ (fsm_output[4])) | (fsm_output[1]) | (fsm_output[7]);
  assign mux_267_nl = MUX_s_1_2_2(mux_tmp_33, or_tmp_23, fsm_output[3]);
  assign mux_266_nl = MUX_s_1_2_2(and_485_cse, (fsm_output[4]), fsm_output[3]);
  assign mux_268_nl = MUX_s_1_2_2(mux_267_nl, mux_266_nl, fsm_output[1]);
  assign mux_265_nl = MUX_s_1_2_2(mux_tmp_264, mux_tmp_263, fsm_output[1]);
  assign mux_269_nl = MUX_s_1_2_2(mux_268_nl, mux_265_nl, fsm_output[2]);
  assign mux_270_nl = MUX_s_1_2_2(mux_269_nl, or_tmp_298, fsm_output[0]);
  assign ecb1_nor_5_seb = ~(mux_270_nl | or_404_cse);
  assign ecb1_or_10_cse = and_307_ssc | and_308_ssc | and_309_ssc | and_310_ssc |
      and_318_ssc | (and_dcpl_279 & and_dcpl_291) | and_320_ssc | and_321_ssc;
  assign ecb1_nor_1_cse = ~(and_305_ssc | and_dcpl_263 | and_dcpl_264 | and_311_ssc
      | and_313_ssc | and_dcpl_277 | and_dcpl_278);
  assign mux_277_nl = MUX_s_1_2_2(mux_37_cse, mux_tmp_273, fsm_output[2]);
  assign mux_275_nl = MUX_s_1_2_2(mux_37_cse, mux_tmp_264, fsm_output[1]);
  assign mux_276_nl = MUX_s_1_2_2(mux_275_nl, mux_tmp_273, fsm_output[2]);
  assign mux_278_nl = MUX_s_1_2_2(mux_277_nl, mux_276_nl, fsm_output[0]);
  assign ecb1_nor_4_seb = ~(mux_278_nl | or_404_cse);
  assign and_301_seb = and_dcpl_257 & and_dcpl_288;
  assign and_560_cse = (fsm_output[2:1]==2'b11);
  assign nor_280_cse = ~((fsm_output[6]) | (fsm_output[1]));
  assign or_349_nl = (fsm_output[3]) | mux_tmp_33;
  assign mux_280_nl = MUX_s_1_2_2(mux_35_cse, or_349_nl, and_560_cse);
  assign mux_281_nl = MUX_s_1_2_2(mux_280_nl, or_tmp_298, fsm_output[0]);
  assign and_322_ssc = (~ mux_281_nl) & and_dcpl_19;
  assign and_323_ssc = and_dcpl_262 & and_dcpl_272;
  assign and_326_ssc = (~ mux_282_itm) & nor_280_cse & and_dcpl_77;
  assign and_329_ssc = (~ mux_282_itm) & (~ (fsm_output[6])) & (fsm_output[1]) &
      and_dcpl_77;
  assign nor_59_cse = ~((fsm_output[4]) | (~ (fsm_output[1])));
  assign or_363_cse = (~ (fsm_output[1])) | (~ (fsm_output[6])) | (fsm_output[7]);
  assign or_358_cse = (~ (fsm_output[4])) | (~ (fsm_output[6])) | (fsm_output[7]);
  assign mux_294_cse = MUX_s_1_2_2(mux_tmp_293, or_572_cse, fsm_output[1]);
  assign nor_286_cse = ~((fsm_output[2:1]!=2'b00));
  assign or_404_cse = (fsm_output[7:6]!=2'b00);
  assign or_409_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[6]);
  assign mux_336_nl = MUX_s_1_2_2(or_572_cse, or_tmp_314, fsm_output[2]);
  assign mux_337_nl = MUX_s_1_2_2(or_409_nl, mux_336_nl, fsm_output[1]);
  assign or_408_nl = and_560_cse | (fsm_output[7:6]!=2'b01);
  assign mux_338_nl = MUX_s_1_2_2(mux_337_nl, or_408_nl, fsm_output[5]);
  assign mux_334_nl = MUX_s_1_2_2(or_tmp_314, mux_tmp_330, fsm_output[2]);
  assign mux_333_nl = MUX_s_1_2_2(or_404_cse, or_572_cse, fsm_output[2]);
  assign or_405_nl = (fsm_output[1]) | mux_333_nl;
  assign mux_335_nl = MUX_s_1_2_2(mux_334_nl, or_405_nl, fsm_output[5]);
  assign mux_339_nl = MUX_s_1_2_2(mux_338_nl, mux_335_nl, fsm_output[4]);
  assign mux_331_nl = MUX_s_1_2_2(mux_tmp_330, or_572_cse, and_560_cse);
  assign or_403_nl = (fsm_output[5]) | mux_331_nl;
  assign or_401_nl = (~((fsm_output[2:1]!=2'b10))) | (fsm_output[7:6]!=2'b01);
  assign or_399_nl = nor_286_cse | (fsm_output[7:6]!=2'b01);
  assign mux_329_nl = MUX_s_1_2_2(or_401_nl, or_399_nl, fsm_output[5]);
  assign mux_332_nl = MUX_s_1_2_2(or_403_nl, mux_329_nl, fsm_output[4]);
  assign mux_340_nl = MUX_s_1_2_2(mux_339_nl, mux_332_nl, fsm_output[3]);
  assign or_396_nl = (fsm_output[5]) | (fsm_output[2]) | (fsm_output[7]) | (~ (fsm_output[6]));
  assign nor_287_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (~ (fsm_output[6])));
  assign nor_288_nl = ~((fsm_output[2]) | (fsm_output[7]) | (~ (fsm_output[6])));
  assign mux_326_nl = MUX_s_1_2_2(nor_287_nl, nor_288_nl, fsm_output[1]);
  assign nand_31_nl = ~((fsm_output[5]) & mux_326_nl);
  assign mux_327_nl = MUX_s_1_2_2(or_396_nl, nand_31_nl, fsm_output[4]);
  assign or_390_nl = (fsm_output[4]) | (~ (fsm_output[5])) | (~ (fsm_output[1]))
      | (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[6]);
  assign mux_328_nl = MUX_s_1_2_2(mux_327_nl, or_390_nl, fsm_output[3]);
  assign mux_341_seb = MUX_s_1_2_2(mux_340_nl, mux_328_nl, fsm_output[0]);
  assign cpkey_or_15_cse = and_393_ssc | and_395_ssc | and_397_ssc | and_398_ssc
      | and_416_ssc | and_418_ssc | and_420_ssc | and_422_ssc;
  assign cpkey_nor_18_cse = ~(and_388_ssc | and_dcpl_324 | and_dcpl_327 | and_400_ssc
      | and_405_ssc | and_dcpl_344 | and_dcpl_346);
  assign mux_365_nl = MUX_s_1_2_2(or_572_cse, mux_tmp_293, fsm_output[1]);
  assign mux_364_nl = MUX_s_1_2_2(or_572_cse, or_tmp_314, fsm_output[1]);
  assign mux_366_nl = MUX_s_1_2_2(mux_365_nl, mux_364_nl, fsm_output[0]);
  assign mux_367_nl = MUX_s_1_2_2(mux_366_nl, mux_tmp_293, fsm_output[4]);
  assign or_442_nl = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[6]) | (~ (fsm_output[7]));
  assign mux_363_nl = MUX_s_1_2_2(mux_294_cse, or_442_nl, fsm_output[4]);
  assign mux_368_nl = MUX_s_1_2_2(mux_367_nl, mux_363_nl, fsm_output[3]);
  assign nor_293_nl = ~(nor_280_cse | (fsm_output[7]));
  assign nor_294_nl = ~((~((~ (fsm_output[1])) | (fsm_output[6]))) | (fsm_output[7]));
  assign mux_361_nl = MUX_s_1_2_2(nor_293_nl, nor_294_nl, fsm_output[0]);
  assign nand_32_nl = ~((fsm_output[4]) & mux_361_nl);
  assign mux_362_nl = MUX_s_1_2_2(or_572_cse, nand_32_nl, fsm_output[3]);
  assign mux_369_nl = MUX_s_1_2_2(mux_368_nl, mux_362_nl, fsm_output[5]);
  assign mux_357_nl = MUX_s_1_2_2(or_tmp_314, mux_tmp_293, fsm_output[1]);
  assign mux_358_nl = MUX_s_1_2_2(mux_357_nl, mux_294_cse, fsm_output[4]);
  assign mux_354_nl = MUX_s_1_2_2(or_572_cse, or_tmp_314, nor_59_cse);
  assign mux_359_nl = MUX_s_1_2_2(mux_358_nl, mux_354_nl, fsm_output[3]);
  assign or_434_nl = (fsm_output[0]) | (~ (fsm_output[1])) | (~ (fsm_output[6]))
      | (fsm_output[7]);
  assign or_433_nl = (fsm_output[0]) | (fsm_output[1]) | (~ (fsm_output[6])) | (fsm_output[7]);
  assign mux_352_nl = MUX_s_1_2_2(or_434_nl, or_433_nl, fsm_output[4]);
  assign or_431_nl = (~((fsm_output[0]) | (fsm_output[1]) | (fsm_output[6]))) | (fsm_output[7]);
  assign mux_351_nl = MUX_s_1_2_2(or_363_cse, or_431_nl, fsm_output[4]);
  assign mux_353_nl = MUX_s_1_2_2(mux_352_nl, mux_351_nl, fsm_output[3]);
  assign mux_360_nl = MUX_s_1_2_2(mux_359_nl, mux_353_nl, fsm_output[5]);
  assign mux_370_seb = MUX_s_1_2_2(mux_369_nl, mux_360_nl, fsm_output[2]);
  assign mux_349_nl = MUX_s_1_2_2(or_61_cse, or_60_cse, fsm_output[1]);
  assign and_382_seb = (~ mux_349_nl) & (fsm_output[5]) & and_dcpl_368;
  assign or_452_cse = (fsm_output[2]) | (fsm_output[4]) | (~ (fsm_output[6])) | (fsm_output[7]);
  assign nor_297_nl = ~((fsm_output[4:1]!=4'b1000));
  assign and_565_nl = (fsm_output[4:1]==4'b0111);
  assign mux_373_nl = MUX_s_1_2_2(nor_297_nl, and_565_nl, fsm_output[0]);
  assign and_425_ssc = mux_373_nl & and_dcpl_45 & (~ (fsm_output[7]));
  assign nor_301_nl = ~((~(nor_286_cse | (fsm_output[4]))) | (fsm_output[7:6]!=2'b10));
  assign nor_302_nl = ~(and_560_cse | (fsm_output[4]) | (~ (fsm_output[6])) | (fsm_output[7]));
  assign mux_377_nl = MUX_s_1_2_2(nor_301_nl, nor_302_nl, fsm_output[5]);
  assign nor_303_nl = ~(((~((fsm_output[2:1]==2'b11))) & (fsm_output[4])) | (fsm_output[7:6]!=2'b01));
  assign nor_304_nl = ~(nor_286_cse | (~ (fsm_output[4])) | (~ (fsm_output[6])) |
      (fsm_output[7]));
  assign mux_376_nl = MUX_s_1_2_2(nor_303_nl, nor_304_nl, fsm_output[5]);
  assign mux_378_nl = MUX_s_1_2_2(mux_377_nl, mux_376_nl, fsm_output[3]);
  assign nand_106_nl = ~((fsm_output[2]) & (fsm_output[4]) & (fsm_output[6]) & (~
      (fsm_output[7])));
  assign or_450_nl = (fsm_output[2]) | (~ (fsm_output[4])) | (~ (fsm_output[6]))
      | (fsm_output[7]);
  assign mux_374_nl = MUX_s_1_2_2(nand_106_nl, or_450_nl, fsm_output[1]);
  assign mux_375_nl = MUX_s_1_2_2(or_452_cse, mux_374_nl, fsm_output[5]);
  assign nor_305_nl = ~((fsm_output[3]) | mux_375_nl);
  assign mux_379_ssc = MUX_s_1_2_2(mux_378_nl, nor_305_nl, fsm_output[0]);
  assign and_427_ssc = and_dcpl_323 & and_dcpl_360 & and_dcpl_77;
  assign and_429_ssc = not_tmp_195 & ((fsm_output[3]) ^ (fsm_output[2])) & nor_274_cse;
  assign nand_107_nl = ~((fsm_output[1]) & (fsm_output[3]) & (fsm_output[4]) & (fsm_output[6]));
  assign mux_380_nl = MUX_s_1_2_2(nand_107_nl, or_tmp_414, fsm_output[2]);
  assign mux_381_nl = MUX_s_1_2_2(mux_380_nl, or_tmp_412, fsm_output[7]);
  assign and_430_ssc = (~ mux_381_nl) & nor_274_cse;
  assign or_92_cse = (~ (fsm_output[5])) | (fsm_output[7]);
  assign nor_308_cse = ~((fsm_output[0]) | (fsm_output[3]));
  assign and_498_cse = sub_1_equal_tmp_6 & exit_ecb2_sva;
  assign or_65_nl = (fsm_output[6:4]!=3'b100);
  assign mux_53_nl = MUX_s_1_2_2(or_65_nl, or_64_cse, fsm_output[3]);
  assign mux_414_nl = MUX_s_1_2_2(mux_53_nl, mux_tmp_412, fsm_output[1]);
  assign or_491_nl = (fsm_output[1]) | (fsm_output[3]) | (~ nor_tmp_73);
  assign mux_415_nl = MUX_s_1_2_2(mux_414_nl, or_491_nl, fsm_output[2]);
  assign and_449_ssc = (~ mux_415_nl) & and_dcpl_77;
  assign or_507_nl = (~((fsm_output[1]) | (~ (fsm_output[7])))) | (fsm_output[4]);
  assign mux_421_nl = MUX_s_1_2_2(or_tmp_446, or_507_nl, fsm_output[0]);
  assign nand_33_nl = ~((fsm_output[3]) & (~ mux_421_nl));
  assign or_506_nl = (fsm_output[3]) | (fsm_output[1]) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_422_nl = MUX_s_1_2_2(nand_33_nl, or_506_nl, fsm_output[5]);
  assign mux_420_nl = MUX_s_1_2_2(or_tmp_446, or_337_cse, fsm_output[3]);
  assign or_505_nl = (fsm_output[5]) | mux_420_nl;
  assign mux_423_nl = MUX_s_1_2_2(mux_422_nl, or_505_nl, fsm_output[2]);
  assign or_503_nl = (~ (fsm_output[0])) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_417_nl = MUX_s_1_2_2(or_503_nl, or_337_cse, fsm_output[3]);
  assign or_500_nl = (fsm_output[3]) | (~ (fsm_output[0])) | (~ (fsm_output[1]))
      | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_418_nl = MUX_s_1_2_2(mux_417_nl, or_500_nl, fsm_output[5]);
  assign or_498_nl = (fsm_output[3]) | (fsm_output[1]) | (fsm_output[7]) | (~ (fsm_output[4]));
  assign or_496_nl = (fsm_output[3]) | (~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign mux_416_nl = MUX_s_1_2_2(or_498_nl, or_496_nl, fsm_output[5]);
  assign mux_419_nl = MUX_s_1_2_2(mux_418_nl, mux_416_nl, fsm_output[2]);
  assign mux_424_itm = MUX_s_1_2_2(mux_423_nl, mux_419_nl, fsm_output[6]);
  assign and_452_ssc = and_dcpl_245 & (fsm_output[1]) & (~ (fsm_output[7])) & (fsm_output[0]);
  assign or_519_nl = (fsm_output[1]) | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]);
  assign mux_435_nl = MUX_s_1_2_2(or_tmp_412, or_519_nl, fsm_output[2]);
  assign mux_436_nl = MUX_s_1_2_2(or_tmp_414, mux_435_nl, fsm_output[7]);
  assign and_453_ssc = (~ mux_436_nl) & and_dcpl_399;
  assign and_448_itm = nor_326_cse & and_dcpl_1 & nor_279_cse & or_290_cse;
  assign or_672_cse = (fsm_output[4:3]!=2'b00);
  assign sub_1_nor_6_cse = ~((aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[2:0]!=3'b000));
  assign and_579_cse = (fsm_output[0]) & (fsm_output[5]);
  assign mux_37_cse = MUX_s_1_2_2(or_tmp_25, and_485_cse, fsm_output[3]);
  assign cpkey_nor_6_cse = ~((z_out_1[2:0]!=3'b000));
  assign nor_326_cse = ~((fsm_output[6:5]!=2'b00));
  assign mux_468_nl = MUX_s_1_2_2(nor_326_cse, (fsm_output[5]), fsm_output[4]);
  assign and_587_nl = sub_1_equal_tmp_6 & exit_ecb2_sva & (fsm_output[0]);
  assign mux_469_nl = MUX_s_1_2_2(mux_tmp_465, mux_468_nl, and_587_nl);
  assign mux_470_nl = MUX_s_1_2_2(mux_469_nl, nor_tmp_73, fsm_output[3]);
  assign mux_466_nl = MUX_s_1_2_2(mux_tmp_465, nor_tmp_73, fsm_output[0]);
  assign mux_467_nl = MUX_s_1_2_2(mux_466_nl, nor_tmp, fsm_output[3]);
  assign mux_471_nl = MUX_s_1_2_2(mux_470_nl, mux_467_nl, fsm_output[1]);
  assign and_588_nl = or_672_cse & (fsm_output[6:5]==2'b11);
  assign mux_472_nl = MUX_s_1_2_2(mux_471_nl, and_588_nl, fsm_output[2]);
  assign or_547_rgt = mux_472_nl | (fsm_output[7]);
  assign and_463_rgt = nor_tmp & and_dcpl_261 & and_dcpl_260;
  assign or_548_cse = (fsm_output[1]) | (fsm_output[3]);
  assign ecb2_or_2_cse = and_dcpl_432 | and_dcpl_451;
  assign or_562_cse = (fsm_output[3]) | (fsm_output[6]);
  assign or_572_cse = (fsm_output[7:6]!=2'b01);
  assign and_593_cse = (fsm_output[7]) & (fsm_output[5]);
  assign or_64_cse = (fsm_output[6:4]!=3'b000);
  assign or_60_cse = (fsm_output[4]) | (~ (fsm_output[6]));
  assign or_61_cse = (~ (fsm_output[4])) | (fsm_output[6]);
  assign mux_51_cse = MUX_s_1_2_2(or_61_cse, or_60_cse, fsm_output[3]);
  assign aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_addr_mx0w1 = MUX_v_8_16_2((buf_rsci_din[7:0]),
      (buf_rsci_din[15:8]), (buf_rsci_din[23:16]), (buf_rsci_din[31:24]), (buf_rsci_din[39:32]),
      (buf_rsci_din[47:40]), (buf_rsci_din[55:48]), (buf_rsci_din[63:56]), (buf_rsci_din[71:64]),
      (buf_rsci_din[79:72]), (buf_rsci_din[87:80]), (buf_rsci_din[95:88]), (buf_rsci_din[103:96]),
      (buf_rsci_din[111:104]), (buf_rsci_din[119:112]), (buf_rsci_din[127:120]),
      z_out_1[3:0]);
  assign ctx_deckey_rsci_data_in_d_mx0w4 = addkey_1_mux_itm ^ aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out;
  assign ctx_deckey_rsci_data_in_d_mx0w5_7_5 = aes_expandEncKey_1_asn_itm_1_7_5 ^
      (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[7:5]);
  assign ctx_deckey_rsci_data_in_d_mx0w5_4 = aes_expandEncKey_1_asn_itm_1_4_0_rsp_0
      ^ (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[4]);
  assign ctx_deckey_rsci_data_in_d_mx0w5_3_0 = aes_expandEncKey_1_asn_itm_1_4_0_rsp_1
      ^ (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[3:0]);
  assign ctx_key_rsci_data_in_d_mx0w1 = ctx_key_rsci_data_out_d ^ addkey_1_mux_itm;
  assign aes_expandEncKey_xor_2_mx0w3 = rcon_0_sva ^ rcon_7_1_sva;
  assign aes_expandEncKey_xor_1_itm_mx0w4 = rcon_2_sva ^ rcon_7_1_sva;
  assign aes_expandEncKey_xor_mx0w3 = rcon_3_sva ^ rcon_7_1_sva;
  assign mux_32_cse = MUX_s_1_2_2(or_tmp_23, or_tmp_22, fsm_output[3]);
  assign mux_35_cse = MUX_s_1_2_2(or_tmp_25, or_tmp_23, fsm_output[3]);
  assign nor_147_cse = ~((fsm_output[3:2]!=2'b00));
  assign and_503_cse = (fsm_output[3:2]==2'b11);
  assign ecb2_ecb2_or_tmp = addkey_1_equal_tmp_11 | exit_ecb2_sva;
  assign exp1_exp1_xnor_psp_sva_1 = ~(aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_1 ^
      aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_0);
  assign addkey_equal_tmp_6_mx0w1 = (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1==4'b0110);
  assign sub_nor_16_cse = ~((aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[3:2]!=2'b00));
  assign addkey_equal_tmp_3_mx0w1 = (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[1:0]==2'b11)
      & sub_nor_16_cse;
  assign cpkey_cpkey_xor_1_cmx_sva_1 = addkey_1_mux_itm ^ ctx_enckey_rsci_data_out_d;
  assign rj_xtime_x_sva_1 = aes_mixColumns_a_sva_1 ^ aes_mixColumns_b_sva_1;
  assign rj_xtime_x_1_sva_1 = aes_mixColumns_b_sva_1 ^ aes_mixColumns_c_sva_1;
  assign rj_xtime_x_2_sva_1 = aes_mixColumns_c_sva_1 ^ aes_mixColumns_d_sva_1;
  assign rj_xtime_x_3_sva_1 = aes_mixColumns_d_sva_1 ^ aes_mixColumns_a_sva_1;
  assign mix_mix_xor_7_cmx_7_5_sva_1 = (aes_mixColumns_d_sva_1[7:5]) ^ (aes_mixColumns_e_sva_1[7:5])
      ^ (rj_xtime_x_3_sva_1[6:4]);
  assign mix_mix_xor_1_cmx_0_sva_1 = (aes_mixColumns_a_sva_1[0]) ^ (aes_mixColumns_e_sva_1[0])
      ^ (rj_xtime_x_sva_1[7]);
  assign rj_xtime_3_mux_nl = MUX_v_2_2_2((rj_xtime_x_3_sva_1[3:2]), (~ (rj_xtime_x_3_sva_1[3:2])),
      rj_xtime_x_3_sva_1[7]);
  assign mix_mix_xor_7_cmx_4_3_sva_1 = (aes_mixColumns_d_sva_1[4:3]) ^ (aes_mixColumns_e_sva_1[4:3])
      ^ rj_xtime_3_mux_nl;
  assign rj_xtime_mux_1_nl = MUX_s_1_2_2((rj_xtime_x_sva_1[0]), (~ (rj_xtime_x_sva_1[0])),
      rj_xtime_x_sva_1[7]);
  assign mix_mix_xor_1_cmx_1_sva_1 = (aes_mixColumns_a_sva_1[1]) ^ (aes_mixColumns_e_sva_1[1])
      ^ rj_xtime_mux_1_nl;
  assign mix_mix_xor_7_cmx_2_sva_1 = (aes_mixColumns_d_sva_1[2]) ^ (aes_mixColumns_e_sva_1[2])
      ^ (rj_xtime_x_3_sva_1[1]);
  assign mix_mix_xor_1_cmx_2_sva_1 = (aes_mixColumns_a_sva_1[2]) ^ (aes_mixColumns_e_sva_1[2])
      ^ (rj_xtime_x_sva_1[1]);
  assign rj_xtime_3_mux_1_nl = MUX_s_1_2_2((rj_xtime_x_3_sva_1[0]), (~ (rj_xtime_x_3_sva_1[0])),
      rj_xtime_x_3_sva_1[7]);
  assign mix_mix_xor_7_cmx_1_sva_1 = (aes_mixColumns_d_sva_1[1]) ^ (aes_mixColumns_e_sva_1[1])
      ^ rj_xtime_3_mux_1_nl;
  assign rj_xtime_mux_nl = MUX_v_2_2_2((rj_xtime_x_sva_1[3:2]), (~ (rj_xtime_x_sva_1[3:2])),
      rj_xtime_x_sva_1[7]);
  assign mix_mix_xor_1_cmx_4_3_sva_1 = (aes_mixColumns_a_sva_1[4:3]) ^ (aes_mixColumns_e_sva_1[4:3])
      ^ rj_xtime_mux_nl;
  assign mix_mix_xor_7_cmx_0_sva_1 = (aes_mixColumns_d_sva_1[0]) ^ (aes_mixColumns_e_sva_1[0])
      ^ (rj_xtime_x_3_sva_1[7]);
  assign mix_mix_xor_1_cmx_7_5_sva_1 = (aes_mixColumns_a_sva_1[7:5]) ^ (aes_mixColumns_e_sva_1[7:5])
      ^ (rj_xtime_x_sva_1[6:4]);
  assign mix_mix_xor_5_cmx_7_5_sva_1 = (aes_mixColumns_c_sva_1[7:5]) ^ (aes_mixColumns_e_sva_1[7:5])
      ^ (rj_xtime_x_2_sva_1[6:4]);
  assign mix_mix_xor_3_cmx_0_sva_1 = (aes_mixColumns_b_sva_1[0]) ^ (aes_mixColumns_e_sva_1[0])
      ^ (rj_xtime_x_1_sva_1[7]);
  assign rj_xtime_2_mux_nl = MUX_v_2_2_2((rj_xtime_x_2_sva_1[3:2]), (~ (rj_xtime_x_2_sva_1[3:2])),
      rj_xtime_x_2_sva_1[7]);
  assign mix_mix_xor_5_cmx_4_3_sva_1 = (aes_mixColumns_c_sva_1[4:3]) ^ (aes_mixColumns_e_sva_1[4:3])
      ^ rj_xtime_2_mux_nl;
  assign rj_xtime_1_mux_1_nl = MUX_s_1_2_2((rj_xtime_x_1_sva_1[0]), (~ (rj_xtime_x_1_sva_1[0])),
      rj_xtime_x_1_sva_1[7]);
  assign mix_mix_xor_3_cmx_1_sva_1 = (aes_mixColumns_b_sva_1[1]) ^ (aes_mixColumns_e_sva_1[1])
      ^ rj_xtime_1_mux_1_nl;
  assign mix_mix_xor_5_cmx_2_sva_1 = (aes_mixColumns_c_sva_1[2]) ^ (aes_mixColumns_e_sva_1[2])
      ^ (rj_xtime_x_2_sva_1[1]);
  assign mix_mix_xor_3_cmx_2_sva_1 = (aes_mixColumns_b_sva_1[2]) ^ (aes_mixColumns_e_sva_1[2])
      ^ (rj_xtime_x_1_sva_1[1]);
  assign rj_xtime_2_mux_1_nl = MUX_s_1_2_2((rj_xtime_x_2_sva_1[0]), (~ (rj_xtime_x_2_sva_1[0])),
      rj_xtime_x_2_sva_1[7]);
  assign mix_mix_xor_5_cmx_1_sva_1 = (aes_mixColumns_c_sva_1[1]) ^ (aes_mixColumns_e_sva_1[1])
      ^ rj_xtime_2_mux_1_nl;
  assign rj_xtime_1_mux_nl = MUX_v_2_2_2((rj_xtime_x_1_sva_1[3:2]), (~ (rj_xtime_x_1_sva_1[3:2])),
      rj_xtime_x_1_sva_1[7]);
  assign mix_mix_xor_3_cmx_4_3_sva_1 = (aes_mixColumns_b_sva_1[4:3]) ^ (aes_mixColumns_e_sva_1[4:3])
      ^ rj_xtime_1_mux_nl;
  assign mix_mix_xor_5_cmx_0_sva_1 = (aes_mixColumns_c_sva_1[0]) ^ (aes_mixColumns_e_sva_1[0])
      ^ (rj_xtime_x_2_sva_1[7]);
  assign mix_mix_xor_3_cmx_7_5_sva_1 = (aes_mixColumns_b_sva_1[7:5]) ^ (aes_mixColumns_e_sva_1[7:5])
      ^ (rj_xtime_x_1_sva_1[6:4]);
  assign aes_mixColumns_d_sva_1 = MUX_v_8_4_2((buf_rsci_din[31:24]), (buf_rsci_din[63:56]),
      (buf_rsci_din[95:88]), (buf_rsci_din[127:120]), {aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_0
      , aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_1});
  assign aes_mixColumns_e_sva_1 = aes_mixColumns_a_sva_1 ^ aes_mixColumns_b_sva_1
      ^ aes_mixColumns_c_sva_1 ^ aes_mixColumns_d_sva_1;
  assign aes_mixColumns_a_sva_1 = MUX_v_8_4_2((buf_rsci_din[7:0]), (buf_rsci_din[39:32]),
      (buf_rsci_din[71:64]), (buf_rsci_din[103:96]), {aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_0
      , aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_1});
  assign aes_mixColumns_c_sva_1 = MUX_v_8_4_2((buf_rsci_din[23:16]), (buf_rsci_din[55:48]),
      (buf_rsci_din[87:80]), (buf_rsci_din[119:112]), {aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_0
      , aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_1});
  assign aes_mixColumns_b_sva_1 = MUX_v_8_4_2((buf_rsci_din[15:8]), (buf_rsci_din[47:40]),
      (buf_rsci_din[79:72]), (buf_rsci_din[111:104]), {aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_0
      , aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_1});
  assign sub_nor_26_cse = ~((aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[3:1]!=3'b000));
  assign addkey_equal_tmp_16 = (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[0]) & sub_nor_26_cse;
  assign addkey_equal_tmp_17 = (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1==4'b0010);
  assign addkey_equal_tmp_18 = (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1==4'b1100);
  assign addkey_equal_tmp_19 = (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1==4'b0100);
  assign addkey_equal_tmp_20 = (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1==4'b1010);
  assign addkey_equal_tmp_21 = (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1==4'b0101);
  assign addkey_equal_tmp_22 = (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[3]) & addkey_1_nor_6_itm;
  assign sub_1_or_tmp = addkey_equal_tmp_16 | addkey_equal_tmp_17 | sub_1_equal_tmp_3
      | addkey_equal_tmp_19 | addkey_equal_tmp_21 | sub_1_equal_tmp_6 | addkey_1_equal_tmp_7
      | addkey_equal_tmp_22 | sub_1_equal_tmp_9 | addkey_equal_tmp_20 | addkey_1_equal_tmp_11
      | addkey_equal_tmp_18 | addkey_1_equal_tmp_13 | addkey_1_equal_tmp_14 | addkey_1_equal_tmp_15;
  assign addkey_1_or_tmp = addkey_equal_tmp_16 | addkey_equal_tmp_17 | addkey_equal_tmp_3_mx0w1
      | addkey_equal_tmp_19 | addkey_equal_tmp_21 | addkey_equal_tmp_6_mx0w1 | addkey_1_equal_tmp_7
      | addkey_equal_tmp_22 | ((aes_expandEncKey_1_asn_itm_1_4_0_rsp_1==4'b1001))
      | addkey_equal_tmp_20 | addkey_1_equal_tmp_11 | addkey_equal_tmp_18 | addkey_1_equal_tmp_13
      | addkey_1_equal_tmp_14 | addkey_1_equal_tmp_15;
  assign cpkey_nor_2_cse = ~((aes_addRoundKey_cpy_i_4_0_sva_1_3_0[3:2]!=2'b00));
  assign cpkey_cpkey_and_7_cse = (aes_addRoundKey_cpy_i_4_0_sva_1_3_0[3]) & addkey_1_nor_6_itm;
  assign cpkey_or_tmp = ((aes_addRoundKey_cpy_i_4_0_sva_1_3_0==4'b0001)) | ((aes_addRoundKey_cpy_i_4_0_sva_1_3_0==4'b0010))
      | ((aes_addRoundKey_cpy_i_4_0_sva_1_3_0[1:0]==2'b11) & cpkey_nor_2_cse) | ((aes_addRoundKey_cpy_i_4_0_sva_1_3_0==4'b0100))
      | ((aes_addRoundKey_cpy_i_4_0_sva_1_3_0==4'b0101)) | ((aes_addRoundKey_cpy_i_4_0_sva_1_3_0==4'b0110))
      | addkey_1_equal_tmp_7 | cpkey_cpkey_and_7_cse | sub_1_equal_tmp_9 | ((aes_addRoundKey_cpy_i_4_0_sva_1_3_0==4'b1010))
      | addkey_1_equal_tmp_11 | sub_1_equal_tmp_3 | addkey_1_equal_tmp_13 | addkey_1_equal_tmp_14
      | addkey_1_equal_tmp_15;
  assign and_dcpl_263 = and_dcpl_262 & and_dcpl_260;
  assign and_dcpl_264 = and_dcpl_262 & and_dcpl_251;
  assign or_tmp_298 = (fsm_output[5:2]!=4'b0010);
  assign mux_tmp_263 = MUX_s_1_2_2(mux_tmp_33, or_tmp_25, fsm_output[3]);
  assign mux_tmp_264 = MUX_s_1_2_2(or_tmp_25, mux_tmp_33, fsm_output[3]);
  assign and_dcpl_266 = nor_286_cse & and_dcpl_77;
  assign and_dcpl_267 = (fsm_output[4:3]==2'b10);
  assign and_dcpl_268 = nor_326_cse & and_dcpl_267;
  assign and_dcpl_269 = and_dcpl_268 & and_dcpl_266;
  assign and_dcpl_270 = and_dcpl_268 & and_dcpl_251;
  assign and_dcpl_271 = (fsm_output[2:1]==2'b10);
  assign and_dcpl_272 = and_dcpl_271 & and_dcpl_77;
  assign and_dcpl_273 = and_dcpl_268 & and_dcpl_272;
  assign and_dcpl_275 = and_560_cse & and_dcpl_77;
  assign and_dcpl_277 = and_dcpl_245 & and_dcpl_272;
  assign and_dcpl_278 = and_dcpl_245 & and_dcpl_275;
  assign and_dcpl_279 = and_dcpl_45 & nor_279_cse;
  assign and_dcpl_282 = and_dcpl_279 & and_dcpl_275;
  assign and_dcpl_283 = and_dcpl_45 & and_dcpl_261;
  assign and_dcpl_284 = and_dcpl_283 & and_dcpl_266;
  assign and_dcpl_285 = and_dcpl_283 & and_dcpl_251;
  assign and_dcpl_287 = and_dcpl_257 & and_dcpl_272;
  assign and_dcpl_288 = and_dcpl_271 & and_dcpl_254;
  assign and_dcpl_291 = and_560_cse & and_dcpl_254;
  assign mux_272_nl = MUX_s_1_2_2(and_485_cse, or_tmp_25, fsm_output[3]);
  assign mux_271_nl = MUX_s_1_2_2((fsm_output[4]), (fsm_output[5]), fsm_output[3]);
  assign mux_tmp_273 = MUX_s_1_2_2(mux_272_nl, mux_271_nl, fsm_output[1]);
  assign or_75_nl = (fsm_output[5:3]!=3'b100);
  assign mux_282_itm = MUX_s_1_2_2(or_75_nl, or_73_cse, fsm_output[2]);
  assign and_dcpl_318 = and_dcpl_283 & and_dcpl_291;
  assign mux_tmp_293 = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), fsm_output[6]);
  assign or_tmp_314 = (fsm_output[7:6]!=2'b10);
  assign or_tmp_315 = (aes_addRoundKey_cpy_i_4_0_sva_1_3_0[0]) | (fsm_output[7:6]!=2'b01);
  assign or_tmp_317 = (fsm_output[5]) | (fsm_output[7]);
  assign or_tmp_320 = (~((~ (aes_addRoundKey_cpy_i_4_0_sva_1_3_0[0])) | (fsm_output[5])))
      | (fsm_output[7]);
  assign or_tmp_321 = (~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[7]);
  assign and_dcpl_319 = and_dcpl_45 & and_dcpl_267;
  assign mux_324_nl = MUX_s_1_2_2((~ or_tmp_22), and_485_cse, fsm_output[1]);
  assign and_dcpl_323 = mux_324_nl & (fsm_output[6]);
  assign and_dcpl_324 = and_dcpl_323 & nor_147_cse & and_dcpl_254;
  assign and_dcpl_325 = (fsm_output[6]) & (~ (fsm_output[3]));
  assign nor_231_nl = ~((~ (fsm_output[1])) | (fsm_output[4]) | (fsm_output[5]));
  assign nor_232_nl = ~((fsm_output[1]) | (~ and_485_cse));
  assign not_tmp_189 = MUX_s_1_2_2(nor_231_nl, nor_232_nl, fsm_output[2]);
  assign and_dcpl_327 = not_tmp_189 & and_dcpl_325 & and_dcpl_77;
  assign mux_tmp_330 = MUX_s_1_2_2((~ (fsm_output[6])), (fsm_output[6]), fsm_output[7]);
  assign and_dcpl_330 = (fsm_output[3:2]==2'b10);
  assign and_dcpl_332 = and_dcpl_323 & and_dcpl_330 & and_dcpl_77;
  assign and_dcpl_333 = (fsm_output[6]) & (fsm_output[3]);
  assign and_dcpl_335 = not_tmp_189 & and_dcpl_333 & and_dcpl_77;
  assign and_dcpl_338 = and_dcpl_323 & and_503_cse & and_dcpl_77;
  assign and_531_nl = (fsm_output[2]) & (fsm_output[1]) & (fsm_output[3]) & (fsm_output[6]);
  assign nor_233_nl = ~((fsm_output[2]) | (fsm_output[1]) | (fsm_output[3]) | (fsm_output[6]));
  assign not_tmp_193 = MUX_s_1_2_2(and_531_nl, nor_233_nl, fsm_output[7]);
  assign and_dcpl_341 = (fsm_output[2]) & (~ (fsm_output[0]));
  assign and_dcpl_342 = ~((fsm_output[5]) | (fsm_output[3]));
  assign nor_235_nl = ~((fsm_output[1]) | nand_99_cse);
  assign nor_236_nl = ~((~ (fsm_output[1])) | (fsm_output[4]) | (fsm_output[6]));
  assign not_tmp_195 = MUX_s_1_2_2(nor_235_nl, nor_236_nl, fsm_output[7]);
  assign and_dcpl_344 = not_tmp_195 & and_dcpl_342 & and_dcpl_341;
  assign nor_238_nl = ~((fsm_output[3:1]!=3'b011) | nand_99_cse);
  assign nor_239_nl = ~((fsm_output[2]) | (fsm_output[1]) | (~ (fsm_output[3])) |
      (fsm_output[4]) | (fsm_output[6]));
  assign not_tmp_196 = MUX_s_1_2_2(nor_238_nl, nor_239_nl, fsm_output[7]);
  assign and_dcpl_346 = not_tmp_196 & nor_274_cse;
  assign and_dcpl_347 = ~((fsm_output[2]) | (fsm_output[0]));
  assign and_dcpl_348 = (~ (fsm_output[5])) & (fsm_output[3]);
  assign nor_241_nl = ~((fsm_output[2]) | (~((fsm_output[1]) & (fsm_output[4]) &
      (fsm_output[6]))));
  assign nor_242_nl = ~((~ (fsm_output[2])) | (fsm_output[1]) | (fsm_output[4]) |
      (fsm_output[6]));
  assign not_tmp_198 = MUX_s_1_2_2(nor_241_nl, nor_242_nl, fsm_output[7]);
  assign and_dcpl_353 = (fsm_output[5:4]==2'b01);
  assign and_dcpl_355 = not_tmp_193 & and_dcpl_353 & (~ (fsm_output[0]));
  assign nor_243_nl = ~((fsm_output[1]) | (fsm_output[4]) | (~ nor_tmp));
  assign nor_244_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[4])) | (fsm_output[5])
      | (fsm_output[6]));
  assign not_tmp_199 = MUX_s_1_2_2(nor_243_nl, nor_244_nl, fsm_output[7]);
  assign and_dcpl_357 = not_tmp_199 & nor_147_cse & (~ (fsm_output[0]));
  assign nor_245_nl = ~((fsm_output[2]) | (~ (fsm_output[1])) | (fsm_output[4]) |
      (~ nor_tmp));
  assign nor_246_nl = ~((~ (fsm_output[2])) | (fsm_output[1]) | (~ (fsm_output[4]))
      | (fsm_output[5]) | (fsm_output[6]));
  assign not_tmp_200 = MUX_s_1_2_2(nor_245_nl, nor_246_nl, fsm_output[7]);
  assign and_dcpl_359 = not_tmp_200 & nor_308_cse;
  assign and_dcpl_360 = (fsm_output[3:2]==2'b01);
  assign and_dcpl_366 = and_dcpl_45 & and_487_cse;
  assign and_dcpl_368 = and_503_cse & and_dcpl_254;
  assign nor_248_nl = ~((fsm_output[1]) | (fsm_output[3]) | (~ (fsm_output[6])));
  assign nor_249_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[3])) | (fsm_output[6]));
  assign not_tmp_203 = MUX_s_1_2_2(nor_248_nl, nor_249_nl, fsm_output[2]);
  assign and_dcpl_377 = (fsm_output[7:6]==2'b01);
  assign nor_250_nl = ~((fsm_output[1]) | (~((fsm_output[5:3]==3'b111))));
  assign nor_251_nl = ~((~ (fsm_output[1])) | (fsm_output[3]) | (fsm_output[4]) |
      (fsm_output[5]));
  assign not_tmp_207 = MUX_s_1_2_2(nor_250_nl, nor_251_nl, fsm_output[2]);
  assign and_dcpl_396 = (fsm_output[2]) & (fsm_output[0]);
  assign and_dcpl_399 = (~ (fsm_output[5])) & (fsm_output[0]);
  assign or_tmp_412 = (fsm_output[1]) | (~ (fsm_output[3])) | (fsm_output[4]) | (fsm_output[6]);
  assign or_tmp_414 = (~ (fsm_output[1])) | (fsm_output[3]) | nand_99_cse;
  assign nor_tmp_73 = (fsm_output[6:4]==3'b111);
  assign nor_tmp_74 = (fsm_output[6:3]==4'b1111);
  assign mux_382_nl = MUX_s_1_2_2(and_dcpl_45, nor_tmp, fsm_output[4]);
  assign mux_383_nl = MUX_s_1_2_2(nor_tmp_73, mux_382_nl, fsm_output[3]);
  assign mux_tmp_384 = MUX_s_1_2_2(nor_tmp_74, mux_383_nl, fsm_output[1]);
  assign mux_385_nl = MUX_s_1_2_2((~ or_64_cse), nor_tmp_73, fsm_output[3]);
  assign mux_tmp_386 = MUX_s_1_2_2(mux_385_nl, nor_tmp_74, fsm_output[1]);
  assign mux_388_itm = MUX_s_1_2_2(or_7_cse, or_8_cse, fsm_output[4]);
  assign mux_389_nl = MUX_s_1_2_2((~ mux_388_itm), nor_tmp_73, fsm_output[3]);
  assign mux_390_nl = MUX_s_1_2_2(mux_389_nl, nor_tmp_74, fsm_output[1]);
  assign mux_tmp_391 = MUX_s_1_2_2(mux_390_nl, mux_tmp_384, fsm_output[2]);
  assign mux_387_nl = MUX_s_1_2_2(mux_tmp_386, mux_tmp_384, fsm_output[2]);
  assign mux_392_nl = MUX_s_1_2_2(mux_tmp_391, mux_387_nl, fsm_output[0]);
  assign or_dcpl_50 = mux_392_nl | (fsm_output[7]);
  assign mux_393_nl = MUX_s_1_2_2((~ mux_388_itm), nor_tmp, fsm_output[3]);
  assign mux_394_nl = MUX_s_1_2_2(mux_393_nl, nor_tmp_74, fsm_output[1]);
  assign mux_395_nl = MUX_s_1_2_2(mux_394_nl, mux_tmp_384, fsm_output[2]);
  assign or_469_nl = (~ (fsm_output[0])) | (aes_addRoundKey_cpy_i_4_0_sva_1_3_0[0]);
  assign mux_396_nl = MUX_s_1_2_2(mux_395_nl, mux_tmp_391, or_469_nl);
  assign and_dcpl_419 = ~(mux_396_nl | (fsm_output[7]));
  assign and_dcpl_420 = and_dcpl_319 & and_dcpl_260;
  assign and_dcpl_425 = nor_tmp & (~ (fsm_output[4])) & and_dcpl_58 & (~((fsm_output[2])
      | (aes_addRoundKey_cpy_i_4_0_sva_1_3_0[0]))) & and_dcpl_254;
  assign and_537_nl = or_548_cse & (fsm_output[6:4]==3'b111);
  assign mux_397_nl = MUX_s_1_2_2(mux_tmp_386, and_537_nl, fsm_output[2]);
  assign or_dcpl_56 = mux_397_nl | (fsm_output[7]);
  assign nor_256_nl = ~((aes_addRoundKey_cpy_i_4_0_sva_1_3_0[0]) | (~((fsm_output[0])
      & (fsm_output[6]) & (fsm_output[5]))));
  assign mux_401_nl = MUX_s_1_2_2(nor_326_cse, nor_256_nl, fsm_output[3]);
  assign nor_257_nl = ~((~ (fsm_output[0])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_400_nl = MUX_s_1_2_2(nor_257_nl, nor_tmp, fsm_output[3]);
  assign mux_402_nl = MUX_s_1_2_2(mux_401_nl, mux_400_nl, fsm_output[4]);
  assign mux_403_nl = MUX_s_1_2_2(mux_402_nl, nor_tmp_74, fsm_output[2]);
  assign nor_258_nl = ~((~ (fsm_output[3])) | (fsm_output[0]) | (fsm_output[6]) |
      (~ (fsm_output[5])));
  assign mux_398_nl = MUX_s_1_2_2(nor_258_nl, nor_tmp, fsm_output[4]);
  assign mux_399_nl = MUX_s_1_2_2(nor_tmp_74, mux_398_nl, fsm_output[2]);
  assign mux_404_nl = MUX_s_1_2_2(mux_403_nl, mux_399_nl, fsm_output[1]);
  assign and_dcpl_426 = ~(mux_404_nl | (fsm_output[7]));
  assign and_dcpl_428 = (fsm_output[5:4]==2'b10);
  assign or_666_cse = (fsm_output[4]) | (fsm_output[0]);
  assign nand_94_nl = ~((fsm_output[0]) & (fsm_output[5]));
  assign mux_407_nl = MUX_s_1_2_2((fsm_output[5]), nand_94_nl, fsm_output[4]);
  assign nor_264_nl = ~((fsm_output[6]) | mux_407_nl);
  assign and_542_nl = or_666_cse & (fsm_output[5]);
  assign mux_406_nl = MUX_s_1_2_2(and_542_nl, and_485_cse, aes_addRoundKey_cpy_i_4_0_sva_1_3_0[0]);
  assign and_546_nl = (fsm_output[6]) & mux_406_nl;
  assign mux_408_nl = MUX_s_1_2_2(nor_264_nl, and_546_nl, fsm_output[3]);
  assign mux_409_nl = MUX_s_1_2_2(mux_408_nl, nor_tmp_74, fsm_output[2]);
  assign and_548_nl = ((fsm_output[3:2]!=2'b00)) & (fsm_output[6:4]==3'b111);
  assign mux_410_nl = MUX_s_1_2_2(mux_409_nl, and_548_nl, fsm_output[1]);
  assign and_dcpl_431 = ~(mux_410_nl | (fsm_output[7]));
  assign and_dcpl_432 = and_dcpl_283 & and_dcpl_275;
  assign nor_126_nl = ~((fsm_output[6:5]!=2'b10));
  assign mux_55_nl = MUX_s_1_2_2(nor_126_nl, nor_tmp, fsm_output[4]);
  assign mux_tmp_412 = MUX_s_1_2_2((~ mux_55_nl), or_64_cse, fsm_output[3]);
  assign or_tmp_446 = (~ (fsm_output[1])) | (~ (fsm_output[7])) | (fsm_output[4]);
  assign mux_tmp_426 = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), fsm_output[5]);
  assign mux_tmp_452 = MUX_s_1_2_2(or_404_cse, (fsm_output[7]), and_579_cse);
  assign and_dcpl_445 = and_dcpl_252 & and_dcpl_255;
  assign and_dcpl_446 = ~(mux_111_itm | (fsm_output[0]));
  assign mux_tmp_465 = MUX_s_1_2_2(nor_326_cse, nor_tmp, fsm_output[4]);
  assign mux_476_nl = MUX_s_1_2_2((~ nor_tmp), or_8_cse, fsm_output[4]);
  assign mux_477_nl = MUX_s_1_2_2(or_4_cse, mux_476_nl, fsm_output[3]);
  assign nand_37_nl = ~((fsm_output[1]) & (~ mux_477_nl));
  assign mux_478_nl = MUX_s_1_2_2(nand_37_nl, or_tmp_116, fsm_output[2]);
  assign mux_479_nl = MUX_s_1_2_2(mux_478_nl, or_tmp_114, fsm_output[7]);
  assign and_dcpl_451 = ~(mux_479_nl | (fsm_output[0]));
  assign mux_tmp_491 = MUX_s_1_2_2((~ (fsm_output[6])), (fsm_output[6]), fsm_output[3]);
  assign or_tmp_545 = (fsm_output[5]) | (fsm_output[3]);
  assign or_tmp_559 = (fsm_output[5]) | (~ (fsm_output[3])) | (fsm_output[7]) | (~
      (fsm_output[6]));
  assign or_626_nl = (~ (fsm_output[5])) | (fsm_output[3]) | (fsm_output[7]) | (fsm_output[6]);
  assign mux_tmp_537 = MUX_s_1_2_2(or_626_nl, or_tmp_559, fsm_output[4]);
  assign mux_540_nl = MUX_s_1_2_2(or_572_cse, or_404_cse, fsm_output[3]);
  assign nand_tmp_50 = ~((fsm_output[5]) & (~ mux_540_nl));
  assign or_585_nl = (~ (fsm_output[2])) | (fsm_output[5]) | (~ (fsm_output[3]));
  assign or_583_nl = (fsm_output[7]) | (fsm_output[2]) | (~ (fsm_output[5])) | (fsm_output[3]);
  assign mux_509_nl = MUX_s_1_2_2(or_585_nl, or_583_nl, fsm_output[1]);
  assign nor_332_nl = ~((fsm_output[4]) | mux_509_nl);
  assign nor_333_nl = ~((fsm_output[1]) | (fsm_output[7]) | (~ (fsm_output[2])) |
      (fsm_output[5]) | (fsm_output[3]));
  assign or_580_nl = (fsm_output[5]) | (~ (fsm_output[3]));
  assign or_579_nl = (~ (fsm_output[5])) | (fsm_output[3]);
  assign mux_507_nl = MUX_s_1_2_2(or_580_nl, or_579_nl, fsm_output[2]);
  assign nor_334_nl = ~((~ (fsm_output[1])) | (fsm_output[7]) | mux_507_nl);
  assign mux_508_nl = MUX_s_1_2_2(nor_333_nl, nor_334_nl, fsm_output[4]);
  assign mux_510_nl = MUX_s_1_2_2(nor_332_nl, mux_508_nl, fsm_output[6]);
  assign aes_expandEncKey_1_i_1_4_2_sva_1_0_mx0c0 = mux_510_nl & (fsm_output[0]);
  assign and_592_nl = (fsm_output[2:1]==2'b11) & (~ mux_51_cse);
  assign nor_335_nl = ~((fsm_output[2]) | (fsm_output[1]) | (fsm_output[3]) | (fsm_output[4])
      | (fsm_output[6]));
  assign mux_511_nl = MUX_s_1_2_2(and_592_nl, nor_335_nl, fsm_output[7]);
  assign aes_expandEncKey_1_i_1_4_2_sva_1_0_mx0c1 = mux_511_nl & and_dcpl_399;
  assign or_2_nl = (fsm_output[4]) | (~ nor_tmp);
  assign or_589_nl = (fsm_output[6:4]!=3'b010);
  assign mux_512_nl = MUX_s_1_2_2(or_2_nl, or_589_nl, fsm_output[3]);
  assign nor_336_nl = ~((fsm_output[1]) | mux_512_nl);
  assign nor_337_nl = ~((~ (fsm_output[1])) | (fsm_output[3]) | (~ (fsm_output[4]))
      | (fsm_output[5]) | (fsm_output[6]));
  assign mux_513_nl = MUX_s_1_2_2(nor_336_nl, nor_337_nl, fsm_output[7]);
  assign aes_expandEncKey_1_i_1_4_2_sva_1_0_mx0c2 = mux_513_nl & and_dcpl_396;
  assign aes_expandEncKey_1_i_1_4_2_sva_1_0_mx0c3 = and_dcpl_319 & and_dcpl_291;
  assign and_277_ssc = and_dcpl_262 & and_dcpl_255;
  assign and_288_ssc = and_dcpl_268 & and_dcpl_275;
  assign and_292_ssc = and_dcpl_279 & and_dcpl_266;
  assign and_293_ssc = and_dcpl_279 & and_dcpl_251;
  assign and_298_ssc = and_dcpl_283 & and_dcpl_272;
  assign and_302_ssc = and_dcpl_257 & and_dcpl_275;
  assign and_304_ssc = and_dcpl_257 & and_dcpl_291;
  assign and_305_ssc = and_dcpl_262 & and_dcpl_266;
  assign and_306_ssc = and_dcpl_262 & and_dcpl_275;
  assign and_307_ssc = and_dcpl_262 & and_dcpl_291;
  assign and_308_ssc = and_dcpl_268 & and_dcpl_260;
  assign and_309_ssc = and_dcpl_268 & and_dcpl_255;
  assign and_310_ssc = and_dcpl_268 & and_dcpl_288;
  assign and_311_ssc = and_dcpl_245 & and_dcpl_266;
  assign and_312_ssc = and_dcpl_245 & and_dcpl_260;
  assign and_313_ssc = and_dcpl_245 & and_dcpl_251;
  assign and_314_ssc = and_dcpl_245 & and_dcpl_255;
  assign and_315_ssc = and_dcpl_245 & and_dcpl_288;
  assign and_316_ssc = and_dcpl_245 & and_dcpl_291;
  assign and_317_ssc = and_dcpl_279 & and_dcpl_272;
  assign and_318_ssc = and_dcpl_279 & and_dcpl_288;
  assign and_320_ssc = and_dcpl_283 & and_dcpl_260;
  assign and_321_ssc = and_dcpl_283 & and_dcpl_255;
  assign and_341_ssc = not_tmp_189 & and_dcpl_325 & and_dcpl_254;
  assign and_352_ssc = not_tmp_193 & (~(or_tmp_22 | (fsm_output[0])));
  assign and_362_ssc = not_tmp_195 & and_dcpl_348 & and_dcpl_347;
  assign and_364_ssc = not_tmp_198 & and_dcpl_348 & (~ (fsm_output[0]));
  assign and_374_ssc = not_tmp_199 & and_dcpl_360 & (~ (fsm_output[0]));
  assign and_500_nl = (fsm_output[2]) & (fsm_output[1]) & (~ (fsm_output[4])) & (fsm_output[6]);
  assign nor_290_nl = ~((fsm_output[2]) | (fsm_output[1]) | (~ (fsm_output[4])) |
      (fsm_output[6]));
  assign mux_348_nl = MUX_s_1_2_2(and_500_nl, nor_290_nl, fsm_output[0]);
  assign and_377_ssc = mux_348_nl & (fsm_output[5]) & (fsm_output[3]) & (~ (fsm_output[7]));
  assign and_384_ssc = not_tmp_203 & and_485_cse & and_dcpl_77;
  assign and_386_ssc = not_tmp_203 & and_485_cse & and_dcpl_254;
  assign and_388_ssc = and_dcpl_323 & nor_147_cse & and_dcpl_77;
  assign and_391_ssc = not_tmp_207 & and_dcpl_377 & (~ (fsm_output[0]));
  assign and_393_ssc = not_tmp_207 & and_dcpl_377 & (fsm_output[0]);
  assign and_395_ssc = and_dcpl_323 & and_dcpl_330 & and_dcpl_254;
  assign and_397_ssc = not_tmp_189 & and_dcpl_333 & and_dcpl_254;
  assign and_398_ssc = and_dcpl_323 & and_dcpl_368;
  assign and_400_ssc = not_tmp_195 & and_dcpl_342 & and_dcpl_347;
  assign and_403_ssc = not_tmp_195 & and_dcpl_342 & (~ (fsm_output[2])) & (fsm_output[0]);
  assign and_405_ssc = not_tmp_198 & and_dcpl_342 & (~ (fsm_output[0]));
  assign and_407_ssc = not_tmp_198 & and_dcpl_342 & (fsm_output[0]);
  assign and_410_ssc = not_tmp_195 & and_dcpl_342 & and_dcpl_396;
  assign and_412_ssc = not_tmp_196 & and_dcpl_399;
  assign and_414_ssc = not_tmp_195 & and_dcpl_348 & and_dcpl_341;
  assign and_416_ssc = not_tmp_195 & and_dcpl_348 & and_dcpl_396;
  assign and_418_ssc = not_tmp_193 & and_dcpl_353 & (fsm_output[0]);
  assign and_420_ssc = not_tmp_199 & nor_147_cse & (fsm_output[0]);
  assign and_422_ssc = not_tmp_200 & (~ (fsm_output[3])) & (fsm_output[0]);
  assign or_446_nl = (fsm_output[4:1]!=4'b0011) | (~ nor_tmp);
  assign mux_372_nl = MUX_s_1_2_2(or_446_nl, or_tmp_114, fsm_output[7]);
  assign nor_296_ssc = ~(mux_372_nl | (fsm_output[0]));
  assign aes_expandEncKey_1_aes_expandEncKey_1_xor_5_nl = (ctx_key_rsci_data_out_d[7])
      ^ (aes_expandEncKey_1_asn_itm_1_7_5[2]);
  assign aes_expandEncKey_1_aes_expandEncKey_1_xor_33_nl = (ctx_key_rsci_data_out_d[7])
      ^ (aes_expandEncKey_1_asn_itm_1_7_5[2]) ^ rcon_7_1_sva;
  assign ecb1_mux1h_4_nl = MUX1HOT_s_1_6_2((ctx_enckey_rsci_data_out_d[7]), (ctx_key_rsci_data_in_d_mx0w1[7]),
      aes_expandEncKey_1_aes_expandEncKey_1_xor_5_nl, aes_expandEncKey_1_aes_expandEncKey_1_xor_33_nl,
      (ctx_deckey_rsci_data_in_d_mx0w4[7]), (ctx_deckey_rsci_data_in_d_mx0w5_7_5[2]),
      {and_425_ssc , mux_379_ssc , and_dcpl_327 , and_427_ssc , and_429_ssc , and_430_ssc});
  assign aes_expandEncKey_1_aes_expandEncKey_1_xor_39_nl = (ctx_key_rsci_data_out_d[6])
      ^ (aes_expandEncKey_1_asn_itm_1_7_5[1]);
  assign aes_expandEncKey_1_aes_expandEncKey_1_xor_27_nl = (ctx_key_rsci_data_out_d[6])
      ^ (aes_expandEncKey_1_asn_itm_1_7_5[1]) ^ rcon_6_sva;
  assign ecb1_mux1h_8_nl = MUX1HOT_s_1_6_2((ctx_enckey_rsci_data_out_d[6]), (ctx_key_rsci_data_in_d_mx0w1[6]),
      aes_expandEncKey_1_aes_expandEncKey_1_xor_39_nl, aes_expandEncKey_1_aes_expandEncKey_1_xor_27_nl,
      (ctx_deckey_rsci_data_in_d_mx0w4[6]), (ctx_deckey_rsci_data_in_d_mx0w5_7_5[1]),
      {and_425_ssc , mux_379_ssc , and_dcpl_327 , and_427_ssc , and_429_ssc , and_430_ssc});
  assign aes_expandEncKey_1_aes_expandEncKey_1_xor_40_nl = (ctx_key_rsci_data_out_d[5])
      ^ (aes_expandEncKey_1_asn_itm_1_7_5[0]);
  assign aes_expandEncKey_1_aes_expandEncKey_1_xor_37_nl = (ctx_key_rsci_data_out_d[5])
      ^ (aes_expandEncKey_1_asn_itm_1_7_5[0]) ^ rcon_5_sva;
  assign ecb1_mux1h_9_nl = MUX1HOT_s_1_6_2((ctx_enckey_rsci_data_out_d[5]), (ctx_key_rsci_data_in_d_mx0w1[5]),
      aes_expandEncKey_1_aes_expandEncKey_1_xor_40_nl, aes_expandEncKey_1_aes_expandEncKey_1_xor_37_nl,
      (ctx_deckey_rsci_data_in_d_mx0w4[5]), (ctx_deckey_rsci_data_in_d_mx0w5_7_5[0]),
      {and_425_ssc , mux_379_ssc , and_dcpl_327 , and_427_ssc , and_429_ssc , and_430_ssc});
  assign aes_expandEncKey_1_aes_expandEncKey_1_xor_41_nl = (ctx_key_rsci_data_out_d[4])
      ^ aes_expandEncKey_1_asn_itm_1_4_0_rsp_0;
  assign aes_expandEncKey_1_aes_expandEncKey_1_xor_31_nl = (ctx_key_rsci_data_out_d[4])
      ^ aes_expandEncKey_1_asn_itm_1_4_0_rsp_0 ^ rcon_4_sva;
  assign ecb1_mux1h_10_nl = MUX1HOT_s_1_6_2((ctx_enckey_rsci_data_out_d[4]), (ctx_key_rsci_data_in_d_mx0w1[4]),
      aes_expandEncKey_1_aes_expandEncKey_1_xor_41_nl, aes_expandEncKey_1_aes_expandEncKey_1_xor_31_nl,
      (ctx_deckey_rsci_data_in_d_mx0w4[4]), ctx_deckey_rsci_data_in_d_mx0w5_4, {and_425_ssc
      , mux_379_ssc , and_dcpl_327 , and_427_ssc , and_429_ssc , and_430_ssc});
  assign aes_expandEncKey_1_aes_expandEncKey_1_xor_42_nl = (ctx_key_rsci_data_out_d[3])
      ^ (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[3]);
  assign aes_expandEncKey_1_aes_expandEncKey_1_xor_25_nl = (ctx_key_rsci_data_out_d[3])
      ^ (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[3]) ^ rcon_3_sva;
  assign ecb1_mux1h_11_nl = MUX1HOT_s_1_6_2((ctx_enckey_rsci_data_out_d[3]), (ctx_key_rsci_data_in_d_mx0w1[3]),
      aes_expandEncKey_1_aes_expandEncKey_1_xor_42_nl, aes_expandEncKey_1_aes_expandEncKey_1_xor_25_nl,
      (ctx_deckey_rsci_data_in_d_mx0w4[3]), (ctx_deckey_rsci_data_in_d_mx0w5_3_0[3]),
      {and_425_ssc , mux_379_ssc , and_dcpl_327 , and_427_ssc , and_429_ssc , and_430_ssc});
  assign aes_expandEncKey_1_aes_expandEncKey_1_xor_43_nl = (ctx_key_rsci_data_out_d[2])
      ^ (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[2]);
  assign aes_expandEncKey_1_aes_expandEncKey_1_xor_35_nl = (ctx_key_rsci_data_out_d[2])
      ^ (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[2]) ^ rcon_2_sva;
  assign ecb1_mux1h_12_nl = MUX1HOT_s_1_6_2((ctx_enckey_rsci_data_out_d[2]), (ctx_key_rsci_data_in_d_mx0w1[2]),
      aes_expandEncKey_1_aes_expandEncKey_1_xor_43_nl, aes_expandEncKey_1_aes_expandEncKey_1_xor_35_nl,
      (ctx_deckey_rsci_data_in_d_mx0w4[2]), (ctx_deckey_rsci_data_in_d_mx0w5_3_0[2]),
      {and_425_ssc , mux_379_ssc , and_dcpl_327 , and_427_ssc , and_429_ssc , and_430_ssc});
  assign aes_expandEncKey_1_aes_expandEncKey_1_xor_44_nl = (ctx_key_rsci_data_out_d[1])
      ^ (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[1]);
  assign aes_expandEncKey_1_aes_expandEncKey_1_xor_29_nl = (ctx_key_rsci_data_out_d[1])
      ^ (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[1]) ^ rcon_1_sva;
  assign ecb1_mux1h_13_nl = MUX1HOT_s_1_6_2((ctx_enckey_rsci_data_out_d[1]), (ctx_key_rsci_data_in_d_mx0w1[1]),
      aes_expandEncKey_1_aes_expandEncKey_1_xor_44_nl, aes_expandEncKey_1_aes_expandEncKey_1_xor_29_nl,
      (ctx_deckey_rsci_data_in_d_mx0w4[1]), (ctx_deckey_rsci_data_in_d_mx0w5_3_0[1]),
      {and_425_ssc , mux_379_ssc , and_dcpl_327 , and_427_ssc , and_429_ssc , and_430_ssc});
  assign aes_expandEncKey_1_aes_expandEncKey_1_xor_45_nl = (ctx_key_rsci_data_out_d[0])
      ^ (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[0]);
  assign aes_expandEncKey_1_aes_expandEncKey_1_xor_23_nl = (ctx_key_rsci_data_out_d[0])
      ^ (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[0]) ^ rcon_0_sva;
  assign ecb1_mux1h_14_nl = MUX1HOT_s_1_6_2((ctx_enckey_rsci_data_out_d[0]), (ctx_key_rsci_data_in_d_mx0w1[0]),
      aes_expandEncKey_1_aes_expandEncKey_1_xor_45_nl, aes_expandEncKey_1_aes_expandEncKey_1_xor_23_nl,
      (ctx_deckey_rsci_data_in_d_mx0w4[0]), (ctx_deckey_rsci_data_in_d_mx0w5_3_0[0]),
      {and_425_ssc , mux_379_ssc , and_dcpl_327 , and_427_ssc , and_429_ssc , and_430_ssc});
  assign ctx_key_rsci_data_in_d = {ecb1_mux1h_4_nl , ecb1_mux1h_8_nl , ecb1_mux1h_9_nl
      , ecb1_mux1h_10_nl , ecb1_mux1h_11_nl , ecb1_mux1h_12_nl , ecb1_mux1h_13_nl
      , ecb1_mux1h_14_nl};
  assign cpkey_or_26_cse = (and_dcpl_366 & and_dcpl_251) | nor_296_ssc;
  assign cpkey_cpkey_nor_2_nl = ~(nor_296_ssc | and_388_ssc | and_dcpl_324 | and_dcpl_327
      | and_391_ssc | and_393_ssc | and_dcpl_332 | and_395_ssc | and_dcpl_335 | and_397_ssc
      | and_dcpl_338 | and_398_ssc | and_403_ssc | and_407_ssc | and_410_ssc | and_412_ssc
      | mux_370_seb);
  assign cpkey_or_18_nl = and_391_ssc | and_414_ssc;
  assign cpkey_or_20_nl = and_dcpl_332 | and_dcpl_335 | and_dcpl_338;
  assign cpkey_or_7_nl = and_dcpl_355 | and_dcpl_357 | and_dcpl_359;
  assign cpkey_mux1h_163_nl = MUX1HOT_s_1_5_2((z_out_1[3]), exp1_exp1_xnor_psp_sva_1,
      aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_0, exp1_1_exp1_1_xnor_psp_sva, exp2_1_exp2_1_xnor_psp_sva,
      {cpkey_or_26_cse , cpkey_or_18_nl , cpkey_or_15_cse , cpkey_or_20_nl , cpkey_or_7_nl});
  assign cpkey_or_21_nl = (~((~(((cpkey_mux1h_163_nl | and_377_ssc) & cpkey_nor_18_cse)
      | and_384_ssc | and_386_ssc | and_403_ssc | and_407_ssc | and_410_ssc | and_412_ssc))
      | mux_370_seb)) | and_382_seb;
  assign cpkey_or_8_nl = and_391_ssc | and_414_ssc | and_dcpl_355 | and_dcpl_357
      | and_dcpl_359 | and_dcpl_332 | and_dcpl_335 | and_dcpl_338;
  assign cpkey_mux1h_165_nl = MUX1HOT_s_1_3_2((z_out_1[2]), (~ aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_1),
      aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_1, {cpkey_or_26_cse , cpkey_or_8_nl
      , cpkey_or_15_cse});
  assign cpkey_or_22_nl = (~((~(((cpkey_mux1h_165_nl | and_377_ssc) & cpkey_nor_18_cse)
      | and_384_ssc | and_386_ssc | and_403_ssc | and_407_ssc | and_410_ssc | and_412_ssc))
      | mux_370_seb)) | and_382_seb;
  assign cpkey_and_6_nl = (z_out_1[1:0]) & (signext_2_1(~ and_377_ssc)) & (signext_2_1(~
      and_dcpl_338));
  assign nor_356_nl = ~(and_dcpl_469 | and_dcpl_470);
  assign mux1h_nl = MUX1HOT_v_2_3_2(cpkey_and_6_nl, 2'b10, 2'b01, {nor_356_nl , and_dcpl_469
      , and_dcpl_470});
  assign cpkey_nor_23_nl = ~(MUX_v_2_2_2(mux1h_nl, 2'b11, and_391_ssc));
  assign cpkey_or_19_nl = and_400_ssc | and_403_ssc | and_422_ssc | and_dcpl_359;
  assign cpkey_cpkey_nor_3_nl = ~(cpkey_nor_23_nl | ({{1{and_398_ssc}}, and_398_ssc})
      | (signext_2_1(cpkey_or_19_nl)));
  assign cpkey_or_11_nl = and_388_ssc | and_dcpl_346 | and_412_ssc | and_416_ssc
      | and_393_ssc | and_414_ssc;
  assign cpkey_nor_21_nl = ~(MUX_v_2_2_2(cpkey_cpkey_nor_3_nl, 2'b11, cpkey_or_11_nl));
  assign cpkey_cpkey_nor_6_nl = ~(MUX_v_2_2_2(cpkey_nor_21_nl, 2'b11, mux_370_seb));
  assign cpkey_or_23_nl = MUX_v_2_2_2(cpkey_cpkey_nor_6_nl, 2'b11, and_382_seb);
  assign ctx_key_rsci_addr_rd_d = {cpkey_cpkey_nor_2_nl , cpkey_or_21_nl , cpkey_or_22_nl
      , cpkey_or_23_nl};
  assign cpkey_cpkey_nor_1_nl = ~(and_dcpl_318 | and_dcpl_324 | and_dcpl_327 | and_341_ssc
      | and_dcpl_332 | and_dcpl_335 | and_dcpl_338 | and_352_ssc | mux_341_seb);
  assign cpkey_or_13_nl = and_dcpl_332 | and_dcpl_335 | and_dcpl_338 | and_352_ssc
      | and_dcpl_355 | and_dcpl_357 | and_dcpl_359 | and_374_ssc;
  assign cpkey_cpkey_mux_nl = MUX_v_2_2_2((aes_addRoundKey_cpy_i_4_0_sva_1_3_0[3:2]),
      ({aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_0 , aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_1}),
      cpkey_or_13_nl);
  assign cpkey_nor_12_nl = ~(and_dcpl_324 | and_dcpl_327 | and_341_ssc | and_dcpl_344
      | and_dcpl_346 | and_362_ssc | and_364_ssc);
  assign cpkey_nand_nl = ~(MUX_v_2_2_2(2'b00, cpkey_cpkey_mux_nl, cpkey_nor_12_nl));
  assign cpkey_cpkey_nor_7_nl = ~(MUX_v_2_2_2(cpkey_nand_nl, 2'b11, mux_341_seb));
  assign nor_357_nl = ~(or_dcpl_83 | or_dcpl_86);
  assign mux1h_1_nl = MUX1HOT_v_2_3_2((aes_addRoundKey_cpy_i_4_0_sva_1_3_0[1:0]),
      2'b10, 2'b01, {nor_357_nl , or_dcpl_83 , or_dcpl_86});
  assign cpkey_nor_14_nl = ~(and_dcpl_344 | and_374_ssc);
  assign cpkey_and_nl = mux1h_1_nl & (signext_2_1(~ and_352_ssc)) & (signext_2_1(cpkey_nor_14_nl));
  assign cpkey_or_6_nl = and_dcpl_324 | and_364_ssc | and_dcpl_355 | and_dcpl_332;
  assign cpkey_nor_13_nl = ~(MUX_v_2_2_2(cpkey_and_nl, 2'b11, cpkey_or_6_nl));
  assign cpkey_cpkey_nor_8_nl = ~(MUX_v_2_2_2(cpkey_nor_13_nl, 2'b11, mux_341_seb));
  assign ctx_key_rsci_addr_wr_d = {cpkey_cpkey_nor_1_nl , cpkey_cpkey_nor_7_nl ,
      cpkey_cpkey_nor_8_nl};
  assign or_382_nl = (fsm_output[5]) | (~ (fsm_output[7]));
  assign mux_318_cse = MUX_s_1_2_2(or_382_nl, or_92_cse, fsm_output[1]);
  assign or_387_nl = (~((fsm_output[4]) | (fsm_output[1]))) | (fsm_output[5]) | (~
      (fsm_output[7]));
  assign or_384_nl = (fsm_output[1]) | (fsm_output[5]) | (~ (fsm_output[7]));
  assign or_671_nl = (~((aes_expandEncKey_1_asn_itm_1_4_0_rsp_1!=4'b0000) | addkey_1_nor_6_itm))
      | mux_318_cse;
  assign or_380_nl = (fsm_output[1]) | (~ (z_out[2])) | (aes_addRoundKey_cpy_i_4_0_sva_1_3_0[0])
      | (~ (fsm_output[5])) | (fsm_output[7]);
  assign mux_319_nl = MUX_s_1_2_2(or_671_nl, or_380_nl, fsm_output[0]);
  assign mux_320_nl = MUX_s_1_2_2(or_384_nl, mux_319_nl, fsm_output[4]);
  assign mux_321_nl = MUX_s_1_2_2(or_387_nl, mux_320_nl, fsm_output[3]);
  assign or_379_nl = ((fsm_output[4]) & (fsm_output[1])) | (fsm_output[5]) | (~ (fsm_output[7]));
  assign or_377_nl = (~ (fsm_output[1])) | (fsm_output[5]) | (~ (fsm_output[7]));
  assign or_375_nl = nor_272_cse | (aes_addRoundKey_cpy_i_4_0_sva_1_3_0[0]) | (~
      (fsm_output[5])) | (fsm_output[7]);
  assign mux_316_nl = MUX_s_1_2_2(or_377_nl, or_375_nl, fsm_output[4]);
  assign mux_317_nl = MUX_s_1_2_2(or_379_nl, mux_316_nl, fsm_output[3]);
  assign mux_322_nl = MUX_s_1_2_2(mux_321_nl, mux_317_nl, fsm_output[2]);
  assign mux_313_nl = MUX_s_1_2_2(or_tmp_317, or_92_cse, fsm_output[4]);
  assign mux_314_nl = MUX_s_1_2_2(or_tmp_320, mux_313_nl, fsm_output[3]);
  assign or_373_nl = (~ (fsm_output[1])) | (fsm_output[7]);
  assign mux_309_nl = MUX_s_1_2_2(or_tmp_321, or_373_nl, or_288_cse);
  assign mux_310_nl = MUX_s_1_2_2(mux_309_nl, or_tmp_321, fsm_output[0]);
  assign or_368_nl = (aes_addRoundKey_cpy_i_4_0_sva_1_3_0[0]) | (fsm_output[5]) |
      (fsm_output[7]);
  assign mux_308_nl = MUX_s_1_2_2(or_tmp_320, or_368_nl, fsm_output[1]);
  assign mux_311_nl = MUX_s_1_2_2(mux_310_nl, mux_308_nl, fsm_output[4]);
  assign mux_306_nl = MUX_s_1_2_2(or_tmp_317, or_92_cse, fsm_output[1]);
  assign mux_307_nl = MUX_s_1_2_2(mux_306_nl, (fsm_output[7]), fsm_output[4]);
  assign mux_312_nl = MUX_s_1_2_2(mux_311_nl, mux_307_nl, fsm_output[3]);
  assign mux_315_nl = MUX_s_1_2_2(mux_314_nl, mux_312_nl, fsm_output[2]);
  assign ctx_key_rsci_re_d = MUX_s_1_2_2(mux_322_nl, mux_315_nl, fsm_output[6]);
  assign mux_301_nl = MUX_s_1_2_2(or_tmp_314, or_tmp_315, nor_59_cse);
  assign mux_300_nl = MUX_s_1_2_2(mux_tmp_293, or_tmp_315, fsm_output[4]);
  assign mux_302_nl = MUX_s_1_2_2(mux_301_nl, mux_300_nl, fsm_output[3]);
  assign mux_297_nl = MUX_s_1_2_2(or_tmp_315, or_tmp_314, fsm_output[1]);
  assign mux_296_nl = MUX_s_1_2_2(mux_tmp_293, or_tmp_314, aes_addRoundKey_cpy_i_4_0_sva_1_3_0[0]);
  assign mux_298_nl = MUX_s_1_2_2(mux_297_nl, mux_296_nl, fsm_output[4]);
  assign mux_295_nl = MUX_s_1_2_2(mux_294_cse, or_363_cse, fsm_output[4]);
  assign mux_299_nl = MUX_s_1_2_2(mux_298_nl, mux_295_nl, fsm_output[3]);
  assign mux_303_nl = MUX_s_1_2_2(mux_302_nl, mux_299_nl, fsm_output[2]);
  assign or_361_nl = (fsm_output[1]) | (fsm_output[6]) | sub_1_equal_tmp_6 | (fsm_output[7]);
  assign mux_290_nl = MUX_s_1_2_2(or_572_cse, or_361_nl, fsm_output[4]);
  assign nand_102_nl = ~((fsm_output[4]) & (fsm_output[1]) & (fsm_output[6]) & (~
      (fsm_output[7])));
  assign mux_291_nl = MUX_s_1_2_2(mux_290_nl, nand_102_nl, fsm_output[3]);
  assign or_359_nl = nor_59_cse | (fsm_output[7:6]!=2'b01);
  assign mux_289_nl = MUX_s_1_2_2(or_359_nl, or_358_cse, fsm_output[3]);
  assign mux_292_nl = MUX_s_1_2_2(mux_291_nl, mux_289_nl, fsm_output[2]);
  assign mux_304_nl = MUX_s_1_2_2(mux_303_nl, mux_292_nl, fsm_output[5]);
  assign or_357_nl = (fsm_output[4:2]!=3'b000) | (aes_addRoundKey_cpy_i_4_0_sva_1_3_0[0])
      | (fsm_output[7:6]!=2'b01);
  assign or_356_nl = (fsm_output[3]) | (~ (fsm_output[4])) | (~ (fsm_output[1]))
      | (~ (fsm_output[6])) | (fsm_output[7]);
  assign or_355_nl = (~ (fsm_output[4])) | (fsm_output[1]) | (~ (fsm_output[6]))
      | (fsm_output[7]);
  assign or_354_nl = (fsm_output[4]) | (~ (fsm_output[1])) | (fsm_output[6]) | sub_1_equal_tmp_6
      | (fsm_output[7]);
  assign mux_286_nl = MUX_s_1_2_2(or_355_nl, or_354_nl, fsm_output[3]);
  assign mux_287_nl = MUX_s_1_2_2(or_356_nl, mux_286_nl, fsm_output[2]);
  assign mux_288_nl = MUX_s_1_2_2(or_357_nl, mux_287_nl, fsm_output[5]);
  assign ctx_key_rsci_we_d = MUX_s_1_2_2(mux_304_nl, mux_288_nl, fsm_output[0]);
  assign ecb1_mux_1_nl = MUX_v_4_2_2((z_out_1[3:0]), aes_addRoundKey_cpy_i_4_0_sva_1_3_0,
      and_dcpl_318);
  assign aes_expandEncKey_aes_expandEncKey_xor_7_nl = (ctx_deckey_rsci_data_out_d[7])
      ^ (addkey_1_mux_itm[7]);
  assign aes_expandEncKey_aes_expandEncKey_xor_5_nl = (ctx_deckey_rsci_data_out_d[7])
      ^ (aes_expandEncKey_1_asn_itm_1_7_5[2]);
  assign aes_expandEncKey_aes_expandEncKey_xor_22_nl = (ctx_deckey_rsci_data_out_d[7])
      ^ (aes_expandEncKey_1_asn_itm_1_7_5[2]) ^ rcon_7_1_sva;
  assign ecb1_mux1h_3_nl = MUX1HOT_s_1_6_2((k_rsci_data_out_d[7]), aes_expandEncKey_aes_expandEncKey_xor_7_nl,
      aes_expandEncKey_aes_expandEncKey_xor_5_nl, aes_expandEncKey_aes_expandEncKey_xor_22_nl,
      (ctx_deckey_rsci_data_in_d_mx0w4[7]), (ctx_deckey_rsci_data_in_d_mx0w5_7_5[2]),
      {and_dcpl_259 , and_322_ssc , and_dcpl_264 , and_323_ssc , and_326_ssc , and_329_ssc});
  assign aes_expandEncKey_aes_expandEncKey_xor_23_nl = (ctx_deckey_rsci_data_out_d[6])
      ^ (addkey_1_mux_itm[6]);
  assign aes_expandEncKey_aes_expandEncKey_xor_24_nl = (ctx_deckey_rsci_data_out_d[6])
      ^ (aes_expandEncKey_1_asn_itm_1_7_5[1]);
  assign aes_expandEncKey_aes_expandEncKey_xor_20_nl = (ctx_deckey_rsci_data_out_d[6])
      ^ (aes_expandEncKey_1_asn_itm_1_7_5[1]) ^ rcon_6_sva;
  assign ecb1_mux1h_15_nl = MUX1HOT_s_1_6_2((k_rsci_data_out_d[6]), aes_expandEncKey_aes_expandEncKey_xor_23_nl,
      aes_expandEncKey_aes_expandEncKey_xor_24_nl, aes_expandEncKey_aes_expandEncKey_xor_20_nl,
      (ctx_deckey_rsci_data_in_d_mx0w4[6]), (ctx_deckey_rsci_data_in_d_mx0w5_7_5[1]),
      {and_dcpl_259 , and_322_ssc , and_dcpl_264 , and_323_ssc , and_326_ssc , and_329_ssc});
  assign aes_expandEncKey_aes_expandEncKey_xor_25_nl = (ctx_deckey_rsci_data_out_d[5])
      ^ (addkey_1_mux_itm[5]);
  assign aes_expandEncKey_aes_expandEncKey_xor_26_nl = (ctx_deckey_rsci_data_out_d[5])
      ^ (aes_expandEncKey_1_asn_itm_1_7_5[0]);
  assign aes_expandEncKey_aes_expandEncKey_xor_18_nl = (ctx_deckey_rsci_data_out_d[5])
      ^ (aes_expandEncKey_1_asn_itm_1_7_5[0]) ^ rcon_5_sva;
  assign ecb1_mux1h_16_nl = MUX1HOT_s_1_6_2((k_rsci_data_out_d[5]), aes_expandEncKey_aes_expandEncKey_xor_25_nl,
      aes_expandEncKey_aes_expandEncKey_xor_26_nl, aes_expandEncKey_aes_expandEncKey_xor_18_nl,
      (ctx_deckey_rsci_data_in_d_mx0w4[5]), (ctx_deckey_rsci_data_in_d_mx0w5_7_5[0]),
      {and_dcpl_259 , and_322_ssc , and_dcpl_264 , and_323_ssc , and_326_ssc , and_329_ssc});
  assign aes_expandEncKey_aes_expandEncKey_xor_27_nl = (ctx_deckey_rsci_data_out_d[4])
      ^ (addkey_1_mux_itm[4]);
  assign aes_expandEncKey_aes_expandEncKey_xor_28_nl = (ctx_deckey_rsci_data_out_d[4])
      ^ aes_expandEncKey_1_asn_itm_1_4_0_rsp_0;
  assign aes_expandEncKey_aes_expandEncKey_xor_16_nl = (ctx_deckey_rsci_data_out_d[4])
      ^ aes_expandEncKey_1_asn_itm_1_4_0_rsp_0 ^ rcon_4_sva;
  assign ecb1_mux1h_17_nl = MUX1HOT_s_1_6_2((k_rsci_data_out_d[4]), aes_expandEncKey_aes_expandEncKey_xor_27_nl,
      aes_expandEncKey_aes_expandEncKey_xor_28_nl, aes_expandEncKey_aes_expandEncKey_xor_16_nl,
      (ctx_deckey_rsci_data_in_d_mx0w4[4]), ctx_deckey_rsci_data_in_d_mx0w5_4, {and_dcpl_259
      , and_322_ssc , and_dcpl_264 , and_323_ssc , and_326_ssc , and_329_ssc});
  assign aes_expandEncKey_aes_expandEncKey_xor_29_nl = (ctx_deckey_rsci_data_out_d[3])
      ^ (addkey_1_mux_itm[3]);
  assign aes_expandEncKey_aes_expandEncKey_xor_30_nl = (ctx_deckey_rsci_data_out_d[3])
      ^ (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[3]);
  assign aes_expandEncKey_aes_expandEncKey_xor_1_nl = (ctx_deckey_rsci_data_out_d[3])
      ^ (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[3]) ^ rcon_3_sva;
  assign ecb1_mux1h_18_nl = MUX1HOT_s_1_6_2((k_rsci_data_out_d[3]), aes_expandEncKey_aes_expandEncKey_xor_29_nl,
      aes_expandEncKey_aes_expandEncKey_xor_30_nl, aes_expandEncKey_aes_expandEncKey_xor_1_nl,
      (ctx_deckey_rsci_data_in_d_mx0w4[3]), (ctx_deckey_rsci_data_in_d_mx0w5_3_0[3]),
      {and_dcpl_259 , and_322_ssc , and_dcpl_264 , and_323_ssc , and_326_ssc , and_329_ssc});
  assign aes_expandEncKey_aes_expandEncKey_xor_31_nl = (ctx_deckey_rsci_data_out_d[2])
      ^ (addkey_1_mux_itm[2]);
  assign aes_expandEncKey_aes_expandEncKey_xor_32_nl = (ctx_deckey_rsci_data_out_d[2])
      ^ (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[2]);
  assign aes_expandEncKey_aes_expandEncKey_xor_17_nl = (ctx_deckey_rsci_data_out_d[2])
      ^ (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[2]) ^ rcon_2_sva;
  assign ecb1_mux1h_19_nl = MUX1HOT_s_1_6_2((k_rsci_data_out_d[2]), aes_expandEncKey_aes_expandEncKey_xor_31_nl,
      aes_expandEncKey_aes_expandEncKey_xor_32_nl, aes_expandEncKey_aes_expandEncKey_xor_17_nl,
      (ctx_deckey_rsci_data_in_d_mx0w4[2]), (ctx_deckey_rsci_data_in_d_mx0w5_3_0[2]),
      {and_dcpl_259 , and_322_ssc , and_dcpl_264 , and_323_ssc , and_326_ssc , and_329_ssc});
  assign aes_expandEncKey_aes_expandEncKey_xor_33_nl = (ctx_deckey_rsci_data_out_d[1])
      ^ (addkey_1_mux_itm[1]);
  assign aes_expandEncKey_aes_expandEncKey_xor_34_nl = (ctx_deckey_rsci_data_out_d[1])
      ^ (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[1]);
  assign aes_expandEncKey_aes_expandEncKey_xor_19_nl = (ctx_deckey_rsci_data_out_d[1])
      ^ (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[1]) ^ rcon_1_sva;
  assign ecb1_mux1h_20_nl = MUX1HOT_s_1_6_2((k_rsci_data_out_d[1]), aes_expandEncKey_aes_expandEncKey_xor_33_nl,
      aes_expandEncKey_aes_expandEncKey_xor_34_nl, aes_expandEncKey_aes_expandEncKey_xor_19_nl,
      (ctx_deckey_rsci_data_in_d_mx0w4[1]), (ctx_deckey_rsci_data_in_d_mx0w5_3_0[1]),
      {and_dcpl_259 , and_322_ssc , and_dcpl_264 , and_323_ssc , and_326_ssc , and_329_ssc});
  assign aes_expandEncKey_aes_expandEncKey_xor_35_nl = (ctx_deckey_rsci_data_out_d[0])
      ^ (addkey_1_mux_itm[0]);
  assign aes_expandEncKey_aes_expandEncKey_xor_36_nl = (ctx_deckey_rsci_data_out_d[0])
      ^ (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[0]);
  assign aes_expandEncKey_aes_expandEncKey_xor_21_nl = (ctx_deckey_rsci_data_out_d[0])
      ^ (aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[0]) ^ rcon_0_sva;
  assign ecb1_mux1h_21_nl = MUX1HOT_s_1_6_2((k_rsci_data_out_d[0]), aes_expandEncKey_aes_expandEncKey_xor_35_nl,
      aes_expandEncKey_aes_expandEncKey_xor_36_nl, aes_expandEncKey_aes_expandEncKey_xor_21_nl,
      (ctx_deckey_rsci_data_in_d_mx0w4[0]), (ctx_deckey_rsci_data_in_d_mx0w5_3_0[0]),
      {and_dcpl_259 , and_322_ssc , and_dcpl_264 , and_323_ssc , and_326_ssc , and_329_ssc});
  assign ctx_deckey_rsci_data_in_d = {ecb1_mux1h_3_nl , ecb1_mux1h_15_nl , ecb1_mux1h_16_nl
      , ecb1_mux1h_17_nl , ecb1_mux1h_18_nl , ecb1_mux1h_19_nl , ecb1_mux1h_20_nl
      , ecb1_mux1h_21_nl};
  assign ecb1_and_nl = (~(and_305_ssc | and_dcpl_263 | and_dcpl_264 | and_306_ssc
      | and_307_ssc | and_dcpl_269 | and_308_ssc | and_dcpl_270 | and_309_ssc | and_dcpl_273
      | and_310_ssc | and_312_ssc | and_314_ssc | and_315_ssc | and_316_ssc)) & ecb1_nor_4_seb;
  assign ecb1_or_14_nl = and_306_ssc | and_317_ssc;
  assign ecb1_or_16_nl = and_dcpl_269 | and_dcpl_270 | and_dcpl_273;
  assign ecb1_or_2_nl = and_dcpl_282 | and_dcpl_284 | and_dcpl_285;
  assign ecb1_mux1h_2_nl = MUX1HOT_s_1_4_2(exp1_exp1_xnor_psp_sva_1, aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_0,
      exp1_1_exp1_1_xnor_psp_sva, exp2_1_exp2_1_xnor_psp_sva, {ecb1_or_14_nl , ecb1_or_10_cse
      , ecb1_or_16_nl , ecb1_or_2_nl});
  assign ecb1_or_17_nl = (((ecb1_mux1h_2_nl & ecb1_nor_1_cse) | and_dcpl_287 | and_302_ssc
      | and_304_ssc | and_312_ssc | and_314_ssc | and_315_ssc | and_316_ssc) & ecb1_nor_4_seb)
      | and_301_seb;
  assign ecb1_ecb1_mux_nl = MUX_s_1_2_2((~ aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_1),
      aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_1, ecb1_or_10_cse);
  assign ecb1_or_18_nl = (((ecb1_ecb1_mux_nl & ecb1_nor_1_cse) | and_dcpl_287 | and_302_ssc
      | and_304_ssc | and_312_ssc | and_314_ssc | and_315_ssc | and_316_ssc) & ecb1_nor_4_seb)
      | and_301_seb;
  assign or_716_nl = or_dcpl_98 | and_dcpl_264 | and_309_ssc | and_320_ssc | and_314_ssc
      | and_313_ssc | and_304_ssc;
  assign mux_564_nl = MUX_v_2_2_2(2'b01, 2'b10, or_716_nl);
  assign ecb1_nor_7_nl = ~(MUX_v_2_2_2(mux_564_nl, 2'b11, and_dcpl_273));
  assign ecb1_nor_6_nl = ~(MUX_v_2_2_2(ecb1_nor_7_nl, 2'b11, and_306_ssc));
  assign ecb1_or_15_nl = and_dcpl_287 | and_311_ssc | and_312_ssc | and_321_ssc |
      and_dcpl_285;
  assign ecb1_ecb1_nor_nl = ~(ecb1_nor_6_nl | ({{1{and_310_ssc}}, and_310_ssc}) |
      (signext_2_1(ecb1_or_15_nl)));
  assign ecb1_and_6_nl = MUX_v_2_2_2(2'b00, ecb1_ecb1_nor_nl, ecb1_nor_4_seb);
  assign or_722_nl = and_dcpl_278 | and_317_ssc | and_307_ssc | and_318_ssc | and_316_ssc
      | and_305_ssc | and_301_seb;
  assign or_728_nl = MUX_v_2_2_2(ecb1_and_6_nl, 2'b11, or_722_nl);
  assign ctx_deckey_rsci_addr_rd_d = {ecb1_and_nl , ecb1_or_17_nl , ecb1_or_18_nl
      , or_728_nl};
  assign i_and_nl = ((aes_expandEncKey_1_asn_itm_1_4_0_rsp_0 & (~(and_dcpl_263 |
      and_dcpl_264 | and_277_ssc | and_dcpl_269 | and_dcpl_270 | and_dcpl_273 | and_288_ssc)))
      | and_dcpl_277 | and_dcpl_278 | and_292_ssc | and_293_ssc | and_dcpl_282 |
      and_dcpl_284 | and_dcpl_285 | and_298_ssc) & ecb1_nor_5_seb;
  assign i_or_nl = and_dcpl_269 | and_dcpl_270 | and_dcpl_273 | and_288_ssc | and_dcpl_282
      | and_dcpl_284 | and_dcpl_285 | and_298_ssc;
  assign i_i_mux_nl = MUX_v_2_2_2((aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[3:2]),
      ({aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_0 , aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_1}),
      i_or_nl);
  assign i_nor_1_nl = ~(and_dcpl_263 | and_dcpl_264 | and_277_ssc | and_dcpl_277
      | and_dcpl_278 | and_292_ssc | and_293_ssc);
  assign i_and_4_nl = i_i_mux_nl & (signext_2_1(i_nor_1_nl)) & ({{1{ecb1_nor_5_seb}},
      ecb1_nor_5_seb});
  assign nor_359_nl = ~(or_dcpl_108 | or_dcpl_111);
  assign mux1h_3_nl = MUX1HOT_v_2_3_2((aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[1:0]),
      2'b10, 2'b01, {nor_359_nl , or_dcpl_108 , or_dcpl_111});
  assign i_nor_2_nl = ~(and_dcpl_277 | and_298_ssc);
  assign i_and_3_nl = mux1h_3_nl & (signext_2_1(~ and_288_ssc)) & (signext_2_1(i_nor_2_nl));
  assign i_or_3_nl = and_dcpl_263 | and_293_ssc | and_dcpl_282 | and_dcpl_269;
  assign i_or_4_nl = MUX_v_2_2_2(i_and_3_nl, 2'b11, i_or_3_nl);
  assign i_and_5_nl = MUX_v_2_2_2(2'b00, i_or_4_nl, ecb1_nor_5_seb);
  assign ctx_deckey_rsci_addr_wr_d = {i_and_nl , i_and_4_nl , i_and_5_nl};
  assign nor_276_nl = ~((~ (fsm_output[4])) | (fsm_output[7]));
  assign nor_277_nl = ~(exit_ecb2_sva | addkey_1_equal_tmp_11 | (fsm_output[7]));
  assign mux_258_nl = MUX_s_1_2_2(nor_276_nl, nor_277_nl, fsm_output[3]);
  assign or_342_nl = (~ (fsm_output[1])) | addkey_1_equal_tmp_11 | (fsm_output[7]);
  assign mux_253_nl = MUX_s_1_2_2(or_342_nl, or_tmp_291, fsm_output[4]);
  assign or_341_nl = ((fsm_output[1]) & addkey_1_equal_tmp_11) | (fsm_output[7]);
  assign mux_252_nl = MUX_s_1_2_2(or_341_nl, or_tmp_291, fsm_output[4]);
  assign or_340_nl = (z_out_1[2:0]!=3'b000);
  assign mux_254_nl = MUX_s_1_2_2(mux_253_nl, mux_252_nl, or_340_nl);
  assign or_339_nl = addkey_1_equal_tmp_11 | (fsm_output[7]);
  assign mux_251_nl = MUX_s_1_2_2(or_339_nl, or_tmp_291, fsm_output[4]);
  assign mux_255_nl = MUX_s_1_2_2(mux_254_nl, mux_251_nl, fsm_output[0]);
  assign mux_256_nl = MUX_s_1_2_2(mux_255_nl, or_337_cse, exit_ecb2_sva);
  assign or_336_nl = (~ addkey_1_equal_tmp_11) | (fsm_output[7]);
  assign mux_249_nl = MUX_s_1_2_2(nor_26_cse, or_336_nl, fsm_output[4]);
  assign mux_248_nl = MUX_s_1_2_2(nor_26_cse, (fsm_output[7]), fsm_output[4]);
  assign mux_250_nl = MUX_s_1_2_2(mux_249_nl, mux_248_nl, exit_ecb2_sva);
  assign mux_257_nl = MUX_s_1_2_2((~ mux_256_nl), mux_250_nl, fsm_output[3]);
  assign mux_259_nl = MUX_s_1_2_2(mux_258_nl, mux_257_nl, fsm_output[2]);
  assign or_334_nl = (~((fsm_output[4:3]!=2'b01))) | (fsm_output[7]);
  assign or_332_nl = nor_279_cse | (fsm_output[7]);
  assign mux_247_nl = MUX_s_1_2_2(or_334_nl, or_332_nl, fsm_output[2]);
  assign mux_260_nl = MUX_s_1_2_2(mux_259_nl, mux_247_nl, fsm_output[5]);
  assign mux_261_nl = MUX_s_1_2_2(mux_260_nl, (fsm_output[7]), fsm_output[6]);
  assign ctx_deckey_rsci_re_d = ~ mux_261_nl;
  assign mux_240_nl = MUX_s_1_2_2((~ or_tmp_281), or_tmp_281, fsm_output[5]);
  assign mux_241_nl = MUX_s_1_2_2(mux_240_nl, mux_tmp_237, fsm_output[2]);
  assign mux_242_nl = MUX_s_1_2_2(mux_tmp_227, mux_241_nl, fsm_output[3]);
  assign mux_238_nl = MUX_s_1_2_2(mux_tmp_237, and_tmp_11, fsm_output[2]);
  assign mux_235_nl = MUX_s_1_2_2((~ (fsm_output[7])), or_tmp_281, fsm_output[5]);
  assign mux_236_nl = MUX_s_1_2_2(mux_235_nl, and_593_cse, fsm_output[2]);
  assign mux_239_nl = MUX_s_1_2_2(mux_238_nl, mux_236_nl, fsm_output[3]);
  assign mux_243_nl = MUX_s_1_2_2(mux_242_nl, mux_239_nl, fsm_output[1]);
  assign or_330_nl = nor_274_cse | (fsm_output[7]);
  assign mux_233_nl = MUX_s_1_2_2(and_593_cse, or_330_nl, fsm_output[2]);
  assign mux_234_nl = MUX_s_1_2_2(mux_tmp_225, mux_233_nl, fsm_output[3]);
  assign mux_244_nl = MUX_s_1_2_2(mux_243_nl, mux_234_nl, fsm_output[4]);
  assign mux_230_nl = MUX_s_1_2_2(and_593_cse, and_tmp_11, fsm_output[3]);
  assign mux_228_nl = MUX_s_1_2_2(mux_tmp_225, and_tmp_11, fsm_output[2]);
  assign mux_229_nl = MUX_s_1_2_2(mux_228_nl, mux_tmp_227, fsm_output[3]);
  assign mux_231_nl = MUX_s_1_2_2(mux_230_nl, mux_229_nl, fsm_output[1]);

  assign or_560_nl = (fsm_output[3]) | (~ nor_tmp_73);
  assign mux_487_nl = MUX_s_1_2_2(mux_tmp_412, or_560_nl, fsm_output[1]);
  assign mux_486_nl = MUX_s_1_2_2(or_64_cse, or_4_cse, fsm_output[3]);
  assign nand_39_nl = ~((fsm_output[1]) & (~ mux_486_nl));
  assign mux_488_nl = MUX_s_1_2_2(mux_487_nl, nand_39_nl, fsm_output[2]);
  assign and_466_nl = (~ mux_488_nl) & and_dcpl_254;
  assign mux_496_nl = MUX_s_1_2_2(mux_tmp_264, mux_35_cse, fsm_output[1]);
  assign mux_495_nl = MUX_s_1_2_2(mux_tmp_263, mux_32_cse, fsm_output[1]);
  assign mux_497_nl = MUX_s_1_2_2(mux_496_nl, mux_495_nl, fsm_output[2]);
  assign and_468_nl = (~ mux_497_nl) & and_dcpl_19 & (fsm_output[0]);
  assign nand_42_nl = ~((fsm_output[4]) & (~ mux_tmp_293));
  assign or_577_nl = (fsm_output[4]) | mux_tmp_293;
  assign mux_503_nl = MUX_s_1_2_2(or_tmp_314, or_577_nl, fsm_output[2]);
  assign mux_504_nl = MUX_s_1_2_2(nand_42_nl, mux_503_nl, fsm_output[1]);
  assign mux_505_nl = MUX_s_1_2_2(mux_504_nl, or_452_cse, fsm_output[5]);
  assign or_575_nl = (~((fsm_output[2]) | (~ (fsm_output[4])))) | (fsm_output[7:6]!=2'b01);
  assign or_574_nl = (fsm_output[4]) | (~ (fsm_output[6])) | (fsm_output[7]);
  assign mux_498_nl = MUX_s_1_2_2(or_tmp_314, or_572_cse, fsm_output[4]);
  assign mux_499_nl = MUX_s_1_2_2(or_574_nl, mux_498_nl, fsm_output[2]);
  assign mux_500_nl = MUX_s_1_2_2(or_575_nl, mux_499_nl, fsm_output[1]);
  assign mux_501_nl = MUX_s_1_2_2(mux_500_nl, or_358_cse, fsm_output[5]);
  assign mux_506_nl = MUX_s_1_2_2(mux_505_nl, mux_501_nl, fsm_output[3]);
  assign and_469_nl = (~ mux_506_nl) & (fsm_output[0]);
  assign or_749_nl = (fsm_output[2]) | (fsm_output[0]) | mux_tmp_491;
  assign nand_123_nl = ~((fsm_output[1]) & (~ mux_tmp_491));
  assign mux_492_nl = MUX_s_1_2_2(or_749_nl, nand_123_nl, fsm_output[4]);
  assign nor_328_nl = ~((~ (fsm_output[2])) | (fsm_output[0]) | (fsm_output[3]) |
      (~ (fsm_output[6])));
  assign nor_329_nl = ~((fsm_output[2]) | (fsm_output[0]) | (fsm_output[3]) | (~
      (fsm_output[6])));
  assign mux_490_nl = MUX_s_1_2_2(nor_328_nl, nor_329_nl, fsm_output[1]);
  assign nand_124_nl = ~((fsm_output[4]) & mux_490_nl);
  assign mux_493_nl = MUX_s_1_2_2(mux_492_nl, nand_124_nl, fsm_output[5]);
  assign or_563_nl = (~ (fsm_output[3])) | (fsm_output[6]);
  assign mux_489_nl = MUX_s_1_2_2(or_563_nl, or_562_cse, fsm_output[2]);
  assign or_750_nl = (fsm_output[5]) | (fsm_output[4]) | (fsm_output[1]) | mux_489_nl;
  assign or_680_nl = (~ (fsm_output[6])) | (fsm_output[5]) | (~ (fsm_output[3]));
  assign nand_114_nl = ~((fsm_output[5]) & (fsm_output[3]));
  assign mux_525_nl = MUX_s_1_2_2(or_tmp_545, nand_114_nl, fsm_output[6]);
  assign mux_526_nl = MUX_s_1_2_2(or_562_cse, mux_525_nl, or_290_cse);
  assign mux_527_nl = MUX_s_1_2_2(or_680_nl, mux_526_nl, fsm_output[4]);
  assign mux_523_nl = MUX_s_1_2_2((fsm_output[3]), (~ or_tmp_545), fsm_output[6]);
  assign nand_47_nl = ~((fsm_output[1:0]==2'b11) & mux_523_nl);
  assign or_605_nl = (fsm_output[1]) | (~((fsm_output[6]) & (fsm_output[5]) & (fsm_output[3])));
  assign mux_524_nl = MUX_s_1_2_2(nand_47_nl, or_605_nl, fsm_output[4]);
  assign mux_528_nl = MUX_s_1_2_2(mux_527_nl, mux_524_nl, fsm_output[2]);
  assign cpkey_cpkey_nor_nl = ~(addkey_1_nor_6_itm | (aes_addRoundKey_cpy_i_4_0_sva_1_3_0!=4'b0000));
  assign or_682_nl = (~ (fsm_output[1])) | (fsm_output[3]);
  assign or_683_nl = (fsm_output[1]) | (~ (fsm_output[3]));
  assign mux_529_nl = MUX_s_1_2_2(or_682_nl, or_683_nl, fsm_output[2]);
  assign nor_350_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[4])
      | (fsm_output[6]));
  assign nor_142_nl = ~((fsm_output[2]) | mux_51_cse);
  assign mux_532_nl = MUX_s_1_2_2(nor_350_nl, nor_142_nl, fsm_output[0]);
  assign or_631_nl = (fsm_output[3]) | (~ (fsm_output[7])) | (fsm_output[6]);
  assign or_630_nl = (fsm_output[3]) | (fsm_output[7]) | (fsm_output[6]);
  assign mux_542_nl = MUX_s_1_2_2(or_631_nl, or_630_nl, fsm_output[5]);
  assign mux_543_nl = MUX_s_1_2_2(nand_tmp_50, mux_542_nl, fsm_output[4]);
  assign or_628_nl = (fsm_output[5]) | (fsm_output[3]) | (~ (fsm_output[7])) | (fsm_output[6]);
  assign mux_541_nl = MUX_s_1_2_2(nand_tmp_50, or_628_nl, fsm_output[4]);
  assign mux_544_nl = MUX_s_1_2_2(mux_543_nl, mux_541_nl, fsm_output[0]);
  assign nand_49_nl = ~((fsm_output[0]) & (~ mux_tmp_537));
  assign mux_545_nl = MUX_s_1_2_2(mux_544_nl, nand_49_nl, fsm_output[2]);
  assign or_627_nl = (fsm_output[7:3]!=5'b10010);
  assign or_625_nl = (~ (fsm_output[3])) | (~ (fsm_output[7])) | (fsm_output[6]);
  assign mux_535_nl = MUX_s_1_2_2(or_625_nl, or_404_cse, fsm_output[5]);
  assign mux_536_nl = MUX_s_1_2_2(mux_535_nl, or_tmp_559, fsm_output[4]);
  assign mux_538_nl = MUX_s_1_2_2(mux_tmp_537, mux_536_nl, fsm_output[0]);
  assign mux_539_nl = MUX_s_1_2_2(or_627_nl, mux_538_nl, fsm_output[2]);
  assign nor_309_nl = ~((~ (fsm_output[3])) | (~ (fsm_output[5])) | (fsm_output[7]));
  assign nor_310_nl = ~(nor_308_cse | (~ (fsm_output[5])) | (fsm_output[7]));
  assign nor_311_nl = ~((fsm_output[3]) | (~ (fsm_output[5])) | (fsm_output[7]));
  assign mux_432_nl = MUX_s_1_2_2(nor_310_nl, nor_311_nl, fsm_output[1]);
  assign mux_433_nl = MUX_s_1_2_2(nor_309_nl, mux_432_nl, fsm_output[2]);
  assign and_571_nl = (fsm_output[6]) & mux_433_nl;
  assign or_645_nl = (~ (fsm_output[3])) | (fsm_output[5]) | (~ (fsm_output[7]));
  assign mux_428_nl = MUX_s_1_2_2(or_92_cse, mux_tmp_426, fsm_output[3]);
  assign mux_429_nl = MUX_s_1_2_2(or_645_nl, mux_428_nl, fsm_output[0]);
  assign nor_86_nl = ~((fsm_output[0]) | (~ (fsm_output[3])));
  assign mux_427_nl = MUX_s_1_2_2(or_92_cse, mux_tmp_426, nor_86_nl);
  assign mux_430_nl = MUX_s_1_2_2(mux_429_nl, mux_427_nl, fsm_output[1]);
  assign or_510_nl = ((fsm_output[3]) & (fsm_output[0])) | (~ (fsm_output[5])) |
      (fsm_output[7]);
  assign or_509_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[5]) | (~
      (fsm_output[7]));
  assign mux_425_nl = MUX_s_1_2_2(or_510_nl, or_509_nl, fsm_output[1]);
  assign mux_431_nl = MUX_s_1_2_2(mux_430_nl, mux_425_nl, fsm_output[2]);
  assign nor_312_nl = ~((fsm_output[6]) | mux_431_nl);
  assign mux_434_nl = MUX_s_1_2_2(and_571_nl, nor_312_nl, fsm_output[4]);
  assign aes_expandEncKey_1_or_3_nl = and_448_itm | mux_434_nl;
  assign aes_expandEncKey_1_mux1h_14_nl = MUX1HOT_v_4_4_2((z_out_1[3:0]), (aes_expandEncKey_read_rom_sbox_rom_map_1_cmp_data_out[3:0]),
      (ctx_deckey_rsci_data_out_d[3:0]), (ctx_key_rsci_data_out_d[3:0]), {aes_expandEncKey_1_or_3_nl
      , and_449_ssc , and_452_ssc , and_453_ssc});
  assign or_774_nl = nor_308_cse | (~ (fsm_output[2]));
  assign or_773_nl = (~ (fsm_output[0])) | (fsm_output[2]);
  assign mux_597_nl = MUX_s_1_2_2(or_774_nl, or_773_nl, fsm_output[3]);
  assign nor_386_nl = ~((~ (fsm_output[6])) | (fsm_output[1]) | (~ (fsm_output[5]))
      | (fsm_output[7]) | mux_597_nl);
  assign or_770_nl = mux_tmp_426 | (~ (fsm_output[0])) | (fsm_output[2]);
  assign mux_594_nl = MUX_s_1_2_2(or_tmp, or_770_nl, fsm_output[3]);
  assign or_769_nl = (fsm_output[3]) | (~ (fsm_output[0])) | or_92_cse | (fsm_output[2]);
  assign mux_595_nl = MUX_s_1_2_2(mux_594_nl, or_769_nl, nor_163_cse);
  assign nor_385_nl = ~((~ or_92_cse) | (fsm_output[2]));
  assign mux_590_nl = MUX_s_1_2_2(or_tmp_611, nor_385_nl, fsm_output[0]);
  assign mux_591_nl = MUX_s_1_2_2(mux_590_nl, or_tmp, fsm_output[3]);
  assign mux_592_nl = MUX_s_1_2_2(mux_tmp_588, mux_591_nl, fsm_output[7]);
  assign nand_126_nl = ~((fsm_output[7]) & (~ mux_tmp_588));
  assign mux_593_nl = MUX_s_1_2_2(mux_592_nl, nand_126_nl, fsm_output[5]);
  assign mux_596_nl = MUX_s_1_2_2(mux_595_nl, mux_593_nl, fsm_output[1]);
  assign nor_387_nl = ~((fsm_output[6]) | mux_596_nl);
  assign mux_598_nl = MUX_s_1_2_2(nor_386_nl, nor_387_nl, fsm_output[4]);
  assign nor_388_nl = ~(mux_598_nl | (and_448_itm & (~ i_nor_3_seb)));
  assign nor_380_nl = ~((fsm_output[2]) | (fsm_output[4]) | (~ (fsm_output[0])));
  assign mux_584_nl = MUX_s_1_2_2(nor_380_nl, mux_tmp_582, fsm_output[3]);
  assign nor_381_nl = ~((fsm_output[3]) | (~ mux_tmp_582));
  assign mux_585_nl = MUX_s_1_2_2(mux_584_nl, nor_381_nl, fsm_output[6]);
  assign or_760_nl = (~ (fsm_output[4])) | (fsm_output[0]);
  assign mux_580_nl = MUX_s_1_2_2((~ nor_tmp_123), or_760_nl, fsm_output[1]);
  assign or_761_nl = (fsm_output[2]) | mux_580_nl;
  assign or_759_nl = (~ (fsm_output[1])) | (~ (fsm_output[4])) | (fsm_output[0]);
  assign mux_577_nl = MUX_s_1_2_2(mux_tmp, or_666_cse, fsm_output[1]);
  assign mux_578_nl = MUX_s_1_2_2(or_759_nl, mux_577_nl, fsm_output[2]);
  assign mux_576_nl = MUX_s_1_2_2(or_tmp_600, or_666_cse, fsm_output[1]);
  assign or_758_nl = (fsm_output[2]) | mux_576_nl;
  assign mux_579_nl = MUX_s_1_2_2(mux_578_nl, or_758_nl, fsm_output[3]);
  assign mux_581_nl = MUX_s_1_2_2(or_761_nl, mux_579_nl, fsm_output[6]);
  assign mux_586_nl = MUX_s_1_2_2(mux_585_nl, (~ mux_581_nl), fsm_output[5]);
  assign mux_574_nl = MUX_s_1_2_2((~ or_tmp_600), nor_tmp_123, fsm_output[1]);
  assign nand_125_nl = ~((fsm_output[2]) & mux_574_nl);
  assign or_754_nl = (fsm_output[2:1]!=2'b00) | mux_tmp;
  assign mux_575_nl = MUX_s_1_2_2(nand_125_nl, or_754_nl, fsm_output[3]);
  assign nor_382_nl = ~((fsm_output[6:5]!=2'b00) | mux_575_nl);
  assign aes_expandEncKey_1_i_aes_expandEncKey_1_i_mux_nl = MUX_s_1_2_2((z_out[0]),
      (z_out_1[0]), aes_expandEncKey_1_i_1_4_2_sva_1_0_mx0c2);
  assign not_1367_nl = ~ and_614_itm;
  assign ecb3_ecb3_and_1_nl = MUX_v_2_2_2(2'b00, (aes_addRoundKey_cpy_i_4_0_sva_1_3_0[3:2]),
      not_1367_nl);
  assign ecb3_mux_3_nl = MUX_s_1_2_2((aes_addRoundKey_cpy_i_4_0_sva_1_3_0[1]), aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_0,
      and_614_itm);
  assign ecb3_mux_4_nl = MUX_s_1_2_2((aes_addRoundKey_cpy_i_4_0_sva_1_3_0[0]), aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_1,
      and_614_itm);
  assign nl_z_out = ({ecb3_ecb3_and_1_nl , ecb3_mux_3_nl , ecb3_mux_4_nl}) + 4'b0001;
  assign z_out = nl_z_out[3:0];
  assign ecb1_ecb1_or_3_nl = (aes_expandEncKey_1_asn_itm_1_4_0_rsp_0 & (~(and_dcpl_492
      | and_dcpl_496 | and_dcpl_498 | and_dcpl_499))) | and_dcpl_503;
  assign ecb1_mux_4_nl = MUX_s_1_2_2((aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[3]),
      (aes_addRoundKey_cpy_i_4_0_sva_1_3_0[3]), and_dcpl_492);
  assign ecb1_ecb1_or_4_nl = (ecb1_mux_4_nl & (~(and_dcpl_496 | and_dcpl_498))) |
      and_dcpl_503;
  assign ecb1_mux1h_27_nl = MUX1HOT_s_1_4_2((aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[2]),
      (aes_addRoundKey_cpy_i_4_0_sva_1_3_0[2]), (ecb2_mux_26_itm[2]), (z_out[3]),
      {ecb1_or_itm , and_dcpl_492 , and_dcpl_496 , and_dcpl_503});
  assign ecb1_or_23_nl = ecb1_mux1h_27_nl | and_dcpl_498;
  assign ecb1_mux1h_28_nl = MUX1HOT_s_1_5_2((aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[1]),
      (aes_addRoundKey_cpy_i_4_0_sva_1_3_0[1]), (ecb2_mux_26_itm[1]), aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_0,
      (z_out[2]), {ecb1_or_itm , and_dcpl_492 , and_dcpl_496 , and_dcpl_498 , and_dcpl_503});
  assign ecb1_mux1h_29_nl = MUX1HOT_s_1_5_2((aes_expandEncKey_1_asn_itm_1_4_0_rsp_1[0]),
      (aes_addRoundKey_cpy_i_4_0_sva_1_3_0[0]), (ecb2_mux_26_itm[0]), aes_expandEncKey_1_i_1_4_2_sva_1_0_rsp_1,
      (z_out[1]), {ecb1_or_itm , and_dcpl_492 , and_dcpl_496 , and_dcpl_498 , and_dcpl_503});
  assign ecb1_ecb1_or_5_nl = and_dcpl_492 | and_dcpl_496 | and_dcpl_499;
  assign nl_z_out_1 = conv_u2u_5_6({ecb1_ecb1_or_3_nl , ecb1_ecb1_or_4_nl , ecb1_or_23_nl
      , ecb1_mux1h_28_nl , ecb1_mux1h_29_nl}) + conv_s2u_2_6({ecb1_ecb1_or_5_nl ,
      1'b1});
  assign z_out_1 = nl_z_out_1[5:0];

  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_5_2;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [4:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_6_2;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [5:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    MUX1HOT_s_1_6_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_7_2;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [6:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_6_2;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [5:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    MUX1HOT_v_2_6_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_7_2;
    input [1:0] input_6;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [6:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    result = result | (input_6 & {2{sel[6]}});
    MUX1HOT_v_2_7_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_6_2;
    input [2:0] input_5;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [5:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    result = result | (input_4 & {3{sel[4]}});
    result = result | (input_5 & {3{sel[5]}});
    MUX1HOT_v_3_6_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_7_2;
    input [2:0] input_6;
    input [2:0] input_5;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [6:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    result = result | (input_4 & {3{sel[4]}});
    result = result | (input_5 & {3{sel[5]}});
    result = result | (input_6 & {3{sel[6]}});
    MUX1HOT_v_3_7_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction
endmodule
